-- todo: implement this, shift register