--===========================================================================--
--
--  S Y N T H E Z I A B L E    SWTBUG ROM   C O R E
--
--  www.OpenCores.Org - April 2003
--  This core adheres to the GNU public license  
--
-- File name      : cfboot68.vhd
--
-- entity name    : boot_rom
--
-- Purpose        : Implements a 256 x 8 ROM containing the
--                  a boot program for Compact Flash
--                  SWTBUG is assumed to reside at
--                  LBA Address $F478 - $F479 of the Compact Flash
--                  Compact Flash is mapped at $8010
--                  ROM Map Switch at $8030 (clear for RAM)
--                  The idea of using a compact flash Boot ROM
--                  Is to save space in the FPGA rather by booting
--                  the ROM into RAM.
--                  
-- Dependencies   : ieee.Std_Logic_1164
--                  ieee.std_logic_unsigned
--                  ieee.std_logic_arith
--
-- Author         : John E. Kent      
--
--===========================================================================----
--
-- Revision History:
--
-- Date:          Revision         Author
-- 11 Apr 2003    0.1              John Kent
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity boot_rom is
  port (
    cs     : in  std_logic;
    addr   : in  std_logic_vector(7 downto 0);
    data   : out std_logic_vector(7 downto 0)
  );
end entity boot_rom;

architecture basic of boot_rom is
  constant width   : integer := 8;
  constant memsize : integer := 256;

  type rom_array is array(0 to memsize-1) of std_logic_vector(width-1 downto 0);

  constant rom_data : rom_array :=
(
"10001110",
"10100111",
"11111110",
"11001110",
"11111111",
"00011000",
"11011111",
"00000100",
"11001110",
"11111111",
"10111111",
"11011111",
"00000110",
"11001110",
"00010000",
"00000000",
"11011111",
"00001000",
"10111101",
"11111111",
"10110011",
"01111110",
"00010000",
"00000000",
"11001110",
"11000000",
"00000000",
"11011111",
"00000000",
"11000110",
"01111000",
"11010111",
"00000011",
"11001110",
"10000000",
"00010000",
"10001101",
"01111011",
"10000110",
"11100000",
"10100111",
"00000110",
"10001101",
"01110101",
"10000110",
"00000001",
"10100111",
"00000001",
"10000110",
"11101111",
"10100111",
"00000111",
"11001110",
"10000000",
"00010000",
"10001101",
"01101000",
"10000110",
"00000001",
"10100111",
"00000010",
"10010110",
"00000011",
"10100111",
"00000011",
"10000110",
"11110100",
"10100111",
"00000100",
"10000110",
"00000000",
"10100111",
"00000101",
"10000110",
"00100000",
"10100111",
"00000111",
"10001101",
"01010010",
"11000110",
"00000010",
"11010111",
"00000010",
"01011111",
"11001110",
"10000000",
"00010000",
"10100110",
"00000111",
"10000101",
"00001000",
"00100111",
"11111010",
"10100110",
"00000000",
"11011110",
"00000000",
"10100111",
"00000000",
"00001000",
"11011111",
"00000000",
"01011010",
"00100110",
"11101011",
"01111010",
"00000000",
"00000010",
"00100110",
"11100110",
"11010110",
"00000011",
"01011100",
"11010111",
"00000011",
"11000001",
"01111010",
"00100110",
"10111101",
"11001110",
"11000000",
"00000000",
"11011111",
"00000100",
"11001110",
"11000100",
"00000000",
"11011111",
"00000110",
"11001110",
"11100000",
"00000000",
"11011111",
"00001000",
"10001101",
"00101011",
"11001110",
"11000000",
"00000000",
"11011111",
"00000100",
"11001110",
"11000100",
"00000000",
"11011111",
"00000110",
"11001110",
"11111100",
"00000000",
"11011111",
"00001000",
"10001101",
"00011010",
"01111111",
"10000000",
"00110000",
"11111110",
"11111111",
"11111110",
"01101110",
"00000000",
"10100110",
"00000111",
"00101011",
"11111100",
"10100110",
"00000111",
"10000101",
"01000000",
"00100111",
"11110110",
"00111001",
"11011110",
"00001000",
"10100111",
"00000000",
"00001000",
"11011111",
"00001000",
"11011110",
"00000100",
"10100110",
"00000000",
"00001000",
"11011111",
"00000100",
"10011100",
"00000110",
"00100110",
"11101110",
"00111001",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000"
);
begin
   data <= rom_data(conv_integer(addr));
end architecture basic;

