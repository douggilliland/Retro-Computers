��   # 0>3 0 ? > > ?? ( t     >=<>: .   &'	8!= 
 
8 '	 
*.
< 9 	
	 .  2 	6> /5#   '4 '  >( .  
+>(0
>(/.  
 	'?  2&     �
�������	�� ��������
��������	���������
� �����
� ����	��������
������	�����
� �����
����
� ������������
�
� �����
�����	����	��������
������	����������   �������  ��������
��
��
�@��z

�����	     �	 ����� D��  ������
��
��
�
�
���� J
�

��
�� ���� �(�
��  �����(��	   �  �Z
���� ��� f� P� �  �������� (�
�	   ��	 �  �
���	����� ��
�� ��
��
��
  �����
�(����F� ���P������	      �	 ��  ����
�	� ����	�
�	�
�	�
�	������
��(�
���
��	 �  ���7  9? @ � �;P� :�  �  �!�����  � �������
���
�
�F� ���J
� �������
��	�
��
�������      �
      ������ ����  ������  ������� ������������	
 T    �����
�   ��}� � ��  ��  �	�	�����	���	 �  ��  �	��	 �@� ���	�	���  �������
  �	��
�	������@��z

���	��	      �		 ������	��
��
����
��
��	 �X� ��
O��PG� +f�]b(�A]� �
X:���
�
�	�(�
�	��
����	����
���	   �	�	���� �����	�� ��	�����  ��� �����
���� ���	�	�	��	���	 ��
    �	������
�  ��
�
� t;OY�5	��`�  ���
  �W�� ����]�G���	��  �(�
��@��
������������
�	 ���
���� ��
�
��	�
���
��	�����
����
��	����
���
��
�
    �	���	 �!���`��� ��M � [O�r� � G�  ������(��	   ���	     �	 ����
�  �	F�

� J���(������	   ���
����
�	X��������	����	� �	 �  ��	����	�  �	� �����	��
��  ��]��	�	����
� � 1 �y ��;O�          P    ��    P                        &                                                                �� ���(�
� a���
����  E�  ���
��	�
�	� ��D��	�����
�� G�	�����	���(�	�(�
� ������	 ��
����	��	�  ( ��


������
�    �  �� ��	��  �����(�
@��
���
��(�
�����
��
����  ��	���	����  � � j]� ? ��	�O� �	����	����@���		 �(�
���� (�
!�a��
��	      �����	�	  � ��
�	��	�	�
��
� ��
!�� ��
��	P��	�	�
�	�
  ��� �  b�	A8. �(O@ �\� �	�	�	�	��	�
(�
���
�	�
�(�
�� �(�
�� (�
���
������
���
  @�	�����	��
�����

� �`�
(�
���
�
��	��
��	��  �	��	�
���	 �	 H��	 �vT�
� ��O��	 W]8 ;��`Y��  


���
  � (�
����	�H�
  �(�
(�H���	���	��	�  (����	�F� �	��	�
� �	��	�� ��	����  ��	
 �    ���� ����    �      

�
"
,
8
H
W
e
r
�
�
� F   / A 8U� � � @ ��� z
� ? ��`���TL@	����NL_  R��	�L@N R��L_  � � �NT �  �� �� ` 	�� �`��   MT R`N �LlL_  L� � ��	�T ���  	�� �`�VC_  	�� �`R��  &!�
���	\�����	�	����(��	   ��	J� �������	�	    ���	    ������	�	����  �(� !�  �� ���	 �  ���������  �a����^�����O� ��C��c>���f��? ;� �]��������	��	� �  ����		(�
��		(�
`��
���!���	!!!���
��������	����
�(��
��	���
	�
  R `O`���  !���	���:�����u������� (�
������
�����������	
   ����	  �  �
����	��	��	����� ���  �	 ���������  ���``�	�R�O�  m�R��N-�	�N���`N-�	�N� �� 
���*  ���Z�	��O�����	������������	��	   ��� (����
�������	�    ����	�	����(�
�	   �	�	�	��	   �������		 ����	���	�    ������
��	��	������
  �	 �� 
 ]���O�+c �#�H��� ��
 ����
�              ��	��	�
���  ��MA �������� ������	�   ��	�  ����T��  �������J

�  �	��
���
��������	���
����
  	�
�[� z
� �	�	? [��#H��� ��Z���  
  ��������  ��	�!@�

� �	
�
�
 �		
	�  �������  �	��	 ���  �������	�  ����	��
��	�   �����
����
����S���
�	 �	  
S	
�)
S	� 8 �� ��y O;`�������3  ������� ����	���P`    �� �u�
�_ � �  ��'�� �@����
4� �P�� �� �� ���� ��	��
[�� �� �  �� � � �� �   �e
�� �  e
� �  W
� �  H
� �  8
� �  ,
� �  "
� �  
� �  �� ��	� � 