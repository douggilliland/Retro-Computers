--!
--! OpenCores PDP-8 Processor
--!	https://opencores.org/projects/pdp8
--!
--! \brief
--!      PDP-8 implementation for the RETRO-EP4CE15 board
--!
--! \details
--! Additional Comments: Build for RETRO-EP4CE15, using EP4CE15 FPGA
--!		http://land-boards.com/blwiki/index.php?title=RETRO-EP4CE15
--! Front Panel
--!		http://land-boards.com/blwiki/index.php?title=PDP-8_Front_Panel#PDP-8_Front_Panel_Assembly_Sheet
--! Uses bin2mif.py utility to convert the DEC bin file to Altera MIF file
--!	Software at:	https://github.com/douggilliland/Linux-68k/tree/master/pdp8
--! VHDL at:	https://github.com/douggilliland/Retro-Computers/tree/master/PDP-8/PDP8_OpenCores/RETRO-EP4CE15_CYCLONE_IV
--!
--! \file
--!      pdp8_top.vhd
--!
--! \author
--!    Joe Manojlovich - joe.manojlovich (at) gmail (dot) com
--!
--!	Doug Gilliland - adapted to EP4CE15 card
--
--------------------------------------------------------------------
--
--  Copyright (C) 2012 Joe Manojlovich
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- version 2.1 of the License.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE. See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.gnu.org/licenses/lgpl.txt
--
--------------------------------------------------------------------
--
-- Comments are formatted for doxygen
--

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
use ieee.numeric_std;
use work.uart_types.all;                        --! UART Types
use work.dk8e_types.all;                        --! DK8E Types
use work.kc8e_types.all;                        --! KC8E Types
use work.kl8e_types.all;                        --! KL8E Types
use work.rk8e_types.all;                        --! RK8E Types
use work.rk05_types.all;                        --! RK05 Types
use work.ls8e_types.all;                        --! LS8E Types
use work.pr8e_types.all;                        --! PR8E Types
use work.cpu_types.all;                         --! CPU Types
use work.sd_types.all;                          --! SD Types
use work.sdspi_types.all;                       --! SPI Types
use work.oct_7seg;

ENTITY pdp8_top IS
  generic(
    invert_reset : std_logic := '1' -- 0 : not invert, 1 invert
    );
  
  PORT ( 
		CLOCK_50 : IN STD_LOGIC;                                     --! Input clock
		RESET : OUT STD_LOGIC;
		-- 
--		SW : IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (others => 'Z');     --! Toggle switches
		sw			 	: in STD_LOGIC_VECTOR(11 downto 0);
		dispPB		: in std_logic;		-- 12 LEDs display select button

--		KEY : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (others => 'Z');    --! Push buttons
		runLED		: out  STD_LOGIC;		-- RUN
		dispLEDs		: out  STD_LOGIC_VECTOR (11 downto 0) := "000000000000";
		dispPCLED	: out  STD_LOGIC;		-- PC is currently displayed on the 12 LEDs
		dispMALED	: out  STD_LOGIC;		-- MQ value?
		dispMDLED	: out  STD_LOGIC;		-- Indicates that the memory data is currently displayed on the 12 LEDs
		dispACLED	: out  STD_LOGIC;		-- Indicates that the Accumulator is currently displayed on the 12 LEDs

		--		LED : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => 'Z');   --! Output green LEDs

		TTY1_TXD : OUT STD_LOGIC;                                    --! UART send line
		TTY1_RXD : IN STD_LOGIC;                                     --! UART receive line
--		TTY2_TXD : OUT STD_LOGIC;                                    --! UART send line
--		TTY2_RXD : IN STD_LOGIC;                                     --! UART receive line	 
--		LPR_TXD : OUT STD_LOGIC;                                     --! LPR send line
--		LPR_RXD : IN STD_LOGIC;                                      --! LPR receive line
--		LPR_CTS : IN STD_LOGIC;
--		LPR_RTS : OUT STD_LOGIC;
--		PTR_TXD : OUT STD_LOGIC;
--		PTR_RXD : IN STD_LOGIC;
--		PTR_CTS : IN STD_LOGIC;
--		PTR_RTS : OUT STD_LOGIC;
		-- USB_CLK_12MHZ : OUT STD_LOGIC; -- FIXME
--		fpMISO : IN STD_LOGIC;
-- 	Front panel is 7 seg LEDs with SPI-ish interface
--		fpMOSI : OUT STD_LOGIC;
--		fpFS : OUT STD_LOGIC;
--		fpSCLK : OUT STD_LOGIC;

--		swLOCK : IN STD_LOGIC;
--		swCONT : IN STD_LOGIC;
--		swBOOT : IN STD_LOGIC;
--		swEXAM : IN STD_LOGIC;
--		swLDADDR : IN STD_LOGIC;
--		swHALT : IN STD_LOGIC;
--		swLDEXTD : IN STD_LOGIC;
--		swSTEP : IN STD_LOGIC;
--		swDEP : IN STD_LOGIC; 
		--
--		swD0 : IN STD_LOGIC;
--		swD1 : IN STD_LOGIC;
--		swD2 : IN STD_LOGIC;
--		swD3 : IN STD_LOGIC;
--		swD4 : IN STD_LOGIC;
--		swD5 : IN STD_LOGIC;
--		swD6 : IN STD_LOGIC;
--		swD7 : IN STD_LOGIC;
--		swD8 : IN STD_LOGIC;
--		swD9 : IN STD_LOGIC;
--		swD10 : IN STD_LOGIC;
--		swD11 : IN STD_LOGIC;
		--
--		swROT0 : IN STD_LOGIC;
--		swROT1 : IN STD_LOGIC;
--		swROT2 : IN STD_LOGIC;
--		swROT3 : IN STD_LOGIC;
--		swROT4 : IN STD_LOGIC;
--		swROT5 : IN STD_LOGIC;
--		swROT6 : IN STD_LOGIC;
--		swROT7 : IN STD_LOGIC;
		--
		sdCS		: OUT STD_LOGIC; --! SD card chip select
		sdCLK		: OUT STD_LOGIC; --! SD card clock
		sdDI		: OUT STD_LOGIC; --! SD card master out slave in
		sdDO		: IN STD_LOGIC; --! SD card master in slave out
		sdCD		: IN STD_LOGIC;
		-- 
--		swCLEAR : IN STD_LOGIC;
--		swWP : IN STD_LOGIC;
	 
		-- Not using the External SRAM but making sure that it's not active
		sramData		: inout std_logic_vector(7 downto 0) := "ZZZZZZZZ";
		sramAddress	: out std_logic_vector(19 downto 0) := x"00000";
		n_sRamWE		: out std_logic :='1';
		n_sRamCS		: out std_logic :='1';
		n_sRamOE		: out std_logic :='1';

		-- Not using the SD RAM but making sure that it's not active
		n_sdRamCas	: out std_logic := '1';		-- CAS on schematic
		n_sdRamRas	: out std_logic := '1';		-- RAS
		n_sdRamWe	: out std_logic := '1';		-- SDWE
		n_sdRamCe	: out std_logic := '1';		-- SD_NCS0
		sdRamClk		: out std_logic := '1';		-- SDCLK0
		sdRamClkEn	: out std_logic := '1';		-- SDCKE0
		sdRamAddr	: out std_logic_vector(14 downto 0) := "000"&x"000";
		sdRamData	: in std_logic_vector(15 downto 0)
    );
END pdp8_top;

 architecture rtl of pdp8_top is
  signal rk8eSTAT		: rk8eSTAT_t;
  signal swCNTL		: swCNTL_t := (others => '0');                       --! Front Panel Control Switches
  signal swROT			: swROT_t := dispIR;                                  --! Front panel rotator switch
  signal swOPT			: swOPT_t;                                           --! PDP-8 options\
  signal swDATA		: swDATA_t;             --! Front panel switches
  signal LED			: std_logic_vector(7 downto 0);
  signal ledDATA		: data_t;
  --
  signal dig_counter			: std_logic_vector (19 downto 0) := (others => '0');
  signal dispstep 				: std_logic := '0';
  signal dispselcnt				: std_logic_vector (2 downto 0) := "000";
  --
  signal dly			: std_logic := '0';         --! Delay used for reset logic
  signal rst			: std_logic := '0';         --! Internal reset line
  signal int_reset	: std_logic;         --! Initial reset line
  signal rst_out		: std_logic;           --! Reset line output to PDP-8
  
  constant max_count : natural := 24000;
  signal op 			: std_logic;
  
  type display_type is (S0, S1, S2, S3, S4, S5);
  signal state: display_type := S0;   
  signal i 				: integer range 0 to 32 := 0;
  --signal i : std_logic_vector(7 downto 0) := (others => '0');
  signal data7			: std_logic_vector(31 downto 0); -- := X"fa00fa00"; -- (others => '0');
  signal ds2, ds1, ds, dsdb : std_logic := '0';

  

begin

	dispLEDs <= ledDATA;
--    constant dispPC     : swROT_t := "000";                     --! Display PC
--    constant dispAC     : swROT_t := "001";                     --! Display AC
--    constant dispIR     : swROT_t := "010";                     --! Display IR
--    constant dispMA     : swROT_t := "011";                     --! Display MA
--    constant dispMD     : swROT_t := "100";                     --! Display MD
--    constant dispMQ     : swROT_t := "101";                     --! Display MQ
--    constant dispST     : swROT_t := "110";                     --! Display ST
--    constant dispSC     : swROT_t := "111";                     --! Display SC
	dispPCLED <= (not swROT(2)) and (not swROT(1)) and (not swROT(0));	--! Display PC
	dispACLED <= (not swROT(2)) and (not swROT(1)) and (    swROT(0));	--! Display AC
	dispMDLED <= (    swROT(2)) and (not swROT(1)) and (not swROT(0));	--! Display MD
	dispMALED <= (    swROT(2)) and (    swROT(1)) and (    swROT(0));	--! Display MA
	
	swOPT.KE8       <= '1'; 
	swOPT.KM8E      <= '1';
	swOPT.TSD       <= '1';
	swOPT.STARTUP   <= '1'; -- Setting the 'STARTUP' bit will cause the PDP8 to boot
	-- to the address in the switch register

	int_reset <= '0';

	-- 2^18 = 256,000, 50M/250K = 200 mS ticks
	process (CLOCK_50) begin
		if rising_edge(CLOCK_50) then
			dig_counter <= dig_counter+1;
		end if;
	end process;

		-- Debounce for display pushbutton
	process (CLOCK_50, dispPB)
	begin
		if rising_edge(CLOCK_50) then
			if dig_counter(17 downto 0) = 0 then
				ds1		<= dispPB;
				ds			<= ds1;
			end if;
		end if;
	end process;

	-- Edge detect/one-shots for step, loadpc, and deposit switches.
	process (CLOCK_50, ds) begin
		if rising_edge(CLOCK_50) then
			ds2		<= ds;
			dispstep <= ds and not ds2;
	   end if;
	end process;
	
-- Display selection
	process (CLOCK_50) begin 
		if rising_edge(CLOCK_50) then
			if dispstep = '1' then
				swROT <= swROT + 1;
			end if;
		end if;
	end process;

	----------------------------------------------------------------------------
	--  RESET signal generator.
	----------------------------------------------------------------------------
	process(CLOCK_50)
	begin
	 if(rising_edge(CLOCK_50)) then
		dly <= ( not(int_reset) and     dly  and not(rst) )
				 or ( not(int_reset) and not(dly) and     rst  );
		rst <= ( not(int_reset) and not(dly) and not(rst) );
	 end if;
	end process;

	rst_out <= rst xor invert_reset ;

	--
	-- Front Panel Data Switches
	--

	swDATA          <= sw;
	--swDATA          <= o"0023";   
	--swDATA          <= o"7400";   

	 compteur : process(CLOCK_50, rst_out)
		  variable count : natural range 0 to max_count := 0;
	 begin
			if rising_edge(CLOCK_50) then
				if count < max_count/2 then
					 op    <='1';
					 count := count + 1;
				elsif count < max_count then
					 op    <='0';
					 count := count + 1;
				else
					 count := 0;
					 op    <='1';
				end if;
		  end if;
	 end process compteur;   

	----------------------------------------------------------------------------
	-- PDP8 Processor
	---------------------------------------------------------------------------    
	iPDP8 : entity work.ePDP8 (rtl) port map (
	 -- System
	 clk      => CLOCK_50,                   --! 50 MHz Clock
	 rst      => rst_out,                    --! Reset Button
	 -- CPU Configuration
	 swCPU    => swPDP8A,                    --! CPU Configured to emulate PDP8A
	 swOPT    => swOPT,                      --! Enable Options
	 -- Real Time Clock Configuration
	 swRTC    => clkDK8EC2,                  --! RTC 50 Hz interrupt
	 -- TTY1 Interfaces
	 tty1BR   => uartBR9600,                 --! TTY1 is 9600 Baud
	 tty1HS   => uartHSnone,                 --! TTY1 has no flow control
	 tty1CTS  => '1',                        --! TTY1 doesn't need CTS
	 tty1RTS  => open,                       --! TTY1 doesn't need RTS
	 tty1RXD  => TTY1_RXD,                   --! TTY1 RXD (to RS-232 interface)
	 tty1TXD  => TTY1_TXD,                   --! TTY1 TXD (to RS-232 interface)
	 -- TTY2 Interfaces
	 tty2BR   => uartBR9600,                 --! TTY2 is 9600 Baud
	 tty2HS   => uartHSnone,                 --! TTY2 has no flow control
	 tty2CTS  => '1',                        --! TTY2 doesn't need CTS
	 tty2RTS  => open,                       --! TTY2 doesn't need RTS
	 tty2RXD  => '1',                        --! TTY2 RXD (tied off)
	 tty2TXD  => open,                       --! TTY2 TXD (tied off)
	 -- LPR Interface
	 lprBR    => uartBR9600,                 --! LPR is 9600 Baud
	 lprHS    => uartHSnone,                 --! LPR has no flow control
	 lprDTR   => '1',                        --! LPR doesn't need DTR
	 lprDSR   => open,                       --! LPR doesn't need DSR
	 lprRXD   => '1',                        --! LPR RXD (tied off)
	 lprTXD   => open,                       --! LPR TXD (tied off)
	 -- Paper Tape Reader Interface
	 ptrBR    => uartBR9600,                 --! PTR is 9600 Baud
	 ptrHS    => uartHSnone,                 --! PTR has no flow control
	 ptrCTS   => '1',                        --! PTR doesn't need CTS
	 ptrRTS   => open,                       --! PTR doesn't need RTS
	 ptrRXD   => '1',                        --! PTR RXD (tied off)
	 ptrTXD   => open,                       --! PTR TXD (tied off)
	 -- Secure Digital Disk Interface
	 sdCD     => sdCD,                        --! SD Card Detect
	 sdWP     => '0',                        --! SD Write Protect
	 sdMISO   => sdDO,                       --! SD Data In
	 sdMOSI   => sdDI,                       --! SD Data Out
	 sdSCLK   => sdCLK,                      --! SD Clock
	 sdCS     => sdCS,                       --! SD Chip Select
	 -- Status
	 rk8eSTAT => rk8eSTAT,                   --! Disk Status (Ignore)
	 -- Switches and LEDS
	 swROT    => swROT,                      --! Data LEDS display PC
	 swDATA   => swDATA,                     --! RK8E Boot Loader Address
	 swCNTL   => swCNTL,                     --! Switches
	 ledRUN => runLED,                       --! Run LED
	 ledDATA => ledDATA,                        --! Data output register
	 ledADDR => open                         --! Address output register
	 );
	 
end rtl;
