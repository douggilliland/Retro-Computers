���@   �  �� � ȃ @ �` @�$ ??? # ?? # ?#!?=#!?=#$#!? #??!#???!$ ?$?$? $ ?!$="===??$  ??????&??                                                                                                                                                                                                �,�|t|�6��      ��;o F`&6�`�Z�Ñ�ZJrrrr�| �1�3�Z��5� ~}| F��6k   ��� 
	Jj	
F
{"@H��	�6
�6�6D� Z�V� t|zb�l(?Z
�}HD��rD�r�|�J
y�D(ZF���?�0� )
   �o�Q�: ��M u�.���� � ������Ϯ�������Ю��������®���˯̽�����������̠����Ҡ��������Ӡ��Ԡ��������Ġ�����������ٍ����Ġ��Š���Ġ�Ӡ�������Ӡ��Ҡ��Ʊ�ˮ�΍������Ըɮ����������Ӡ��Π�� ���n��l� >A���~��&��J� �    �� n��4��c�F��&��& � � @H1�fn�b�l��y /�   ��& ���F���F ��n6��,��r��{ H�.b愑���{֌�   ��� ���� 2��ޑ����d��6k��\���� ����ݏ ^a�?���^����e�?$�^��?�/a?��!�?�X� ?�o���?$��凿d�Q��� ����3�<�ce�?! �X@���r"    = 8 ��?�Q����h�iQ  �@��!pP�q�� h^���Q�Se�R����z��F�X#$�V��R���6Ѐ5Ј���" "RP �\� ߌ �� �            �@�����o 0����%���                     h�                 #? @ �� ������sR�       ��"��"��"��T+DO�L�6� ��T��A��e�$��RC&�D��Ͱ�����o���� ߌ �� l�_���[�bbh@r#f0&gg[V�� `���� }��``�h'0&aibZ���geY���d\i�a�`d��`�h��40704'#!.0&�?�@F�R����(�b�� �PR��$2F�/~�tn8ri��8pisD��(�D07oiD��� p	88F87"7Sk@     @ e	c�R��f~�%�/Rϐg��.�a6�[V�`���[�V ��`���   #0b7big��Q�6Uigc�\)eT�6Pf��g�a\�d��3�(�4��\��e����h�4�(�Ū��0�l�|X��a�bV���/R �RIQ�:1&� ��(�Ꜧ�(?�3�8`/�4�33CD!7D 4�O�4F376���T��e7�3@b8n4Ui�S�ef�~3�ai6 9Wi����ѫaW��9��Q.�8/~��� `6H"����D��b��� ��c�e5�T�T5�fΚR��U5��)���U�5`/�4����U(�37&�l��͙�)���X�!�A �!8o�|kW��Zb#�]e||��!.q|/Q�aV���/� ��6���/�a���KTa�%R��V����C �6�"����è �2274P)2P)Ԫ�a9����2P)R��V���~TR��T�$R	�T9$T	 & �Ry�UU	�U�$Q	2ae��9SKT��U�Hؾ%  � �  %�/���kta�(?H�t9�T�U��S ���44b33b7bq�����34&3 ?�����9b���R��_b�V���_��R� 629�b ��^����  � 6�9r6�n_�z/)~ ~\)a��ɤ"��"��%�S�x#�� �� �� �� �� �� �R	�@2Ri�7:�j\g�ag�V����� ��|� ���6�. ����ہ��6� ��É�� ���ǉ�� ���4�h�x�x�x�{$"f9�oX�~	tj�6? s3�aY��%��6�?3�������Q��a�p!�#3b!!�1��* ��&(?�!����##���P�2&S�q1�J/��1pn�Ѯ�*1`.�"~�1&3��ę�E"3b&rw&w�z��"Xt�9�j�����t9�p!��X����I%H/3�O3�KaH�� �2Ti24a�4Xi�٪�R�b9��  X���� ��4�/�j�$5bE(/�ȯ�5�G�/��5(/~G��5�33b!4����D� t4(/���SU�$4J
��& � Q	4�jQ2��*���4�PT�$3�3�aY��3�F6�D�*�~��Q�(��Vn���~��mK 5�(/�E�����^��g�ag�6j)� �3Qi4�nQ �5�/~�� F�H�j�&$d��a���:?�  b���6���/�Ϩ����D� �6�"`���`/�ۢ`���@/��`���`/�� ������K��"��&�H/�5�� �6�" ��G@.�5&����   	   R�
" '$"#�%2gf�ke�rf��e�CV �a���r�fB,f�"VՇec�V��V����U"Kv��X(���@/���tN�o � ��H@� /�Ϣ����"6�b�/\�� ��?�(��?�+� �6�"��������É�
.

� �C6&7(/�s�?�	�]�7�)\ϛV �d� 6�`��HA�����4U6 Y������M����橒��vՊs$���������blx#OyUOw��3��3; P�Vi}n_6C"@��?��6����Փk ? #�J9i)�s�9pn#bh�?~���*#�/� ��p��-�[�2�l#�J2 >?��ը`�2c�99@"�#� �q.0�"����e��#�/�7��k7bb�k �,������ ���@ x��ficX���� �-��H �(6�!�慅4cH����/����6��6���R��p9! ��b9b2�b�j�&\)J!.�b��l12s2�D!d�"�(���B�=&aa�a��a_���2�?�C����9&S �7�/f���ad��� 3�!!b00&�3�4r44cba3�!�4' /��!� n3&7�J�D�'��&,Ɖ����-R(���-f��+� ���l�à���,¨����'�.�����D	�
�!��",��(?�&�,�g�.����=��(/������-a.=�(��B/~-������,������>�� � ��\�����
�D	��@@f,�o~76-�b�l���\g��L(?�7�@\)\g�\)��h� = (�����(��� /�����/����E���bnj���2�Οj�cɬR��V>��/�΢2i ߘ p	�ǀ�J�&V���V~���V~�Ղ΂|� ��j��8�6 � $p���� 3R�����  ����)y9� @ ` ��!.�s��G��Z�p�(h�Oj	% .OO}�6�Z3b0W�?��wR��c���R���8 �U��~��pI��ǉ���kpA�%tG��f态&p��P)c��R���&Q�����mkQ���k���lp.��/S�H��s�|H>al�����&�p�/~͒�p�G/~Β݊la � Tk�p��A@�al@ kR��p9�a� !�Z�=ЛR���m��f���                                                                                                                                                                                                    ��V)���? D�„b�&��,V~� /��&��"������ ����t"Pt��S�� .֜b�l�&��&ֻJ�����(����b�a̫��/H �0������/�����* ��b(����&�?ٜ���b!���4��t�֫p(�hO�j%� O�Omk�a�Ol�7~�
�%�/�p��T�$c	�R��<2�Ui(�݄iݑJ�(/~*�!�⨦����q*�~�*�"��h��/Ѳb��&+J.J�����cΚR��pE�(@��~��X��&T.�&�_���c��c��l�نk �B�&������ `��� �Ѡ/�خ�݋l;k;�$&����  Up	�������������/  pP�c��R��� �$'''&/p�%'m����$c'c&c%mk  �QF�n��dn! �i��R)�N�/�N�c�R��o��p�%�J[��Z��Z��\��;

@�ζj@%� ��K� �$piM%bLmkY��hO�]O�O�/�M�L�NLB�L�� ����������Yf   � ����������Q��T��F����Y�@�p�{�~�b����r�ʖD �op�"iD��D����D��D��D��D��D��D�� "$$&m�&#�*~z�vN� "r����N$""Ⱥ���D �ƺ+ ����Z�7a��7�H����@{�8��G���S�g�(�S{�غ�~#� $�j�DyʘD�ID]�҂D֒DڒDޒD�D�D�D�D�D��D��D� ��m��i$��������ƒʒђՒْݒ�DD��D ��/����e�����v��Ph� ��/;�G��x&���owP�G�=w ����:}�Om����f!f��?���� ������ʫ��_�m�� !��U�T�� �� @��%��������� r	���Dm p	����h 	I P�o�������D�$������������D �#�*��[��@���o4������Z� `���`H�g P�D �  /�#F#�+ 	�D� o	Ό�rk��~�$@/@��$Fb#iD�s� �#�Jmp��m�p(��\�%�/j�>�)��?om���� ����ֈ6���/�ʨD� �' $!��D� �$@.Hq� ������&>$&���� ���� �t �6�"  �dh���ֈ� �`��6�"���� �%&f'<b$�k ����aʛ\[�Vw��� $Z֛�5�q���%��~�$�H�6��(/���Q��0������f�fgf    ��̾��S��;�
  :bDs	q$�:(/�= ��$/�#�p��!"�"P.$�"��(q.�&��SE�F�/��Q��" ��#w@ �t�!Cb�$�(��#�/�"�#!.""b#�/��"�/��("�J�]��"�$tn��d�#�#�h��J]����݊ ]	$�K� �(4堾(�k�k; c	�T�$R	�U9���2iI YD 0��� �"Qn#i(�� �/��� �#$B�����  ##&$h/� �$�b�b(fn(�$��q���J�(&"$����\)ā� @!�J!�d�C"\!��\)�� #���F�(#H/!�d"Q ��"��ċ = 
�"Qo�"��!�� �&�&*U/ (�(%b�*bU �((&&�&)U/ (ᰰ�tp~���9i)�@� Q�'bU
�Q'�&U/
Q&%bU
�Q%��Q/� �'D.'&b&�%.%�k @+'"'n*&"&n)%"%�k �(.�6Viz�
�.��\�� �(6�H�,��/�/��R��p��������L� ��Ի�$�F����j ��ә� ��.&�/&�&�+ \	��ˁ_�lp�X.y6ViPL6[)��>�� ����(��FbȀ�D!�=0!/�(��!�!!>`怭B;(���(����&(6)6*6+6� ��a�W��b�����2�*�����V����$6%6&6'6�$�%r&r'r�z    T$��p�@ ��%b nj�U(�� $뻫T$��;���K�E�&�p��a�� m����"PQ�Qe� $$&� �(���) Qo�)b ������!�(�(�'��+b �&�+bU �Ѐ&(�'�&*U/ ��(%B�+bU �((&'�&)U/ ((�iQ'�%�&)U/ %Q&��/!�"�i�a� � % �h� � �/�׋ 'a'�&�!&�%�!%�� �+a.+n*!.*n)!.)�k!(b ��~��<b+bD+�*.*)b���&����+b((&*�''&��� �Q�� Qa��0~��&� ��%�%b(&�('��$�kn �$$&%.�/�خ%�/���0&b\B�g\Ya�!����#�/\ �+&r%� ��Q��(�c�+b�*��ق���&/�%�'&&('&�%�'�&&@/�%��؞%%&�Ƚ ($)b%*b&+b'�k )���%(/&�/�(�!$�(����b@!�!!b>�/���@��H��!�J��K�ƈ���� ��'�@�&�+ ($�/��)%b���j�$�k ��)bH�)�*.*+b+�(�K�� �%H/�%&b&�'.'$d�ػ��ي׋�%�)�/���כ �($�$�(��Ȁ����a���biV��R	 c9I9 I  Њ�*I�^PT�$R	�U9�� PQ%�ȣ��;�[6�jm�RϐT7��9&c��R��92& � J9�*Q7�Q8�R��Q9��B�iD m�e������ $nn�nn��n��� �h%�%mk&�/�'�t�_����a6����R��p���e��9�Kc������D�&                                                                                                                                                                                                 �������?�      L��L�Oj%�i6���F?�$"ei��~e	�,}|{*��% ���        � f{      �        �ꤊ z� � �    � 7   �     � �   _
`F��! ������P�"�oѠ��o/�&� �����  ��mlU�%�`{�H\	�0��tn��b�\�"��ǒҼ6��p �� ���KMɀ� ��~�{�&��BNlN�8Nz0�NtN�8NN4zJ
��

�m� yP�g�, �������'��+�q��!�s��&sK�*!��"��*p'+o',�+ ���f�h������?�??r�>�����H�!�h�N!��w?&@�N�L�_ZXH���N`���_
C���e��aQ�U���HI�H?$��HB?&@���!��x N1�y �H!�ۂ%����H!�ƀ���H!���&�Aۡ(B`�N!�y�$�^���Q�$~#M?S�$Q�/MS�K�i���[#�7?�V�������#9�?ۡ �ad��^��H!� ��a?�i�� ?���� �^��H0!�h���	� ��A���f(��� ���?��?H&�X�N!�x����BN�X���Ӑ?H�!�h�N!���A���f(��񿈑ؿI&�?���� ����/���6��?Cc�����P�� W?��H!�����H0!�o�!xC`�8��(H0?V�H�?�BOK[�b��H0!�o��#?x��_�_��_=}T� ����O�4?`����H���#?C��8`C��8`c#��p( �#�H!�#�T�5?ad(?�?�?Y$�?�d(b[�KB��$� ��u�?F��_�5�?BNf�J�3\����o     �Q-�L�MI�KJ�S����3 ��� ��&ѐ; �	H���� �� �q�☭���&��&��&���܆�
. �T�چ������"��b�!.��b ���H.�l��D� �QL�ѐ��@/��  �A��B�Ҩ����J���M `   �!>�@>H1���b������r��D끲��b��b��c��b�j�2 ���b��&��9      � �� � ������ N���Z��9������� ��V��`/�(�������.
�蒊b���!�����{ �����x��&���!�͙���j�fn��!�蓕&H��@�� �眗&����˃ `� �o��$�H�� ���"��7��9      �h/�!���b��j��"��?���@�(/��J܃�ꢈ��8��J  ��b�(/������Ȣ�V����9��c�(���8H
�!��A��B Ѐ�侢���" FV��q�� !���&�?���A��B�T�� ��� ��������+��" 


��H��"�B� j��h�,�b�	� �Y�Y���`O�E�P�U�R4�VE�R2�V#e K�;	"		" 3GQP��"�+HHBHL"��B�	�	
#�y	%p ���G_`��ͤ����e� U�	���SgcXN_S[NcWS4��3j0��� �Y���`U�		$		D3U�3��3�N�NP��%�W��ԗS����q                                                                                                                                                                                                 � �5TXVC`L �1�4ՒN`�`x�y6y'q.��,����* ���&`��Fw�(w�&�Áǔ�J֮ⷋl�жt���'���                         ��hw�&7�yŁ���Ф� �eߒ�n���� ��&�&�t�B��B�v�.�,u�{�@��8�ހ%�� ���⁢�ڟ���-�&-Ƒ�+k&����!�ʑ�������߃ l��=(��(���(/���-�k��'��'|�w����w��r��w�>�����0��&��)��~��(���+v8�� Η��  �ҁ'��'��'��"�����t������r���|���:[9��/e|6�n�[�B���S�a�                 �����٧�b�폓3�&RiU9$	  �1&��� 	 ` t��7��7�[�	�N��7�@�@߈@�h�����x@�h�@� ߘ@@i�ߨ@�i�@����@ g�@����� ��B�H�g P�����Fj ���4���� ��cA�d��É�A�J��K���VI�1�  F[�/�ʲ���s�(P��F�J�P���/r� ���q�pyuX��Y��� � [��[�kʡft�� ����ʨ��(���[�J��"���Zɀ�� ~��Dԭ���t@�� F���z ��7��K �ʿb��b�ob[�k   �[�������"!��<��p�{U�\�/!.�0b��h�ji7i	��Ѓ � [�\�n"�p��B�j.`�٤:& �h�����FziF6&h���`{P�\��/�&0�&��&t��˨/\v��"����B�z ���)��(��˭ �� ���KUɀ� ��~�{�&��B�l��8�z0��t��8��4zJ
��

��܊ � +  ����K��� ����|u�'s�,׀�E��(}�(���@/}\m�*��/��6�l�r��6��|rq>}�?�m�웊 �줋�-B��t.�'�fI-�&.�&׻6��     \��o נ?�t"���׺B��t��'�F&ӻ�㹌� ���ng �,�


B��h 
��@ `�6�#�c��ǁ����;� �� �� �� �� �� �� Ϧ���:fh~��66���zF���z��q)��}��4�,�7|\���� 5j"�i6�;-&.?b����:&�A�A{�0 ���/j<��i�,�q蘑Oà�t�<��| �����<tt~t�<o�	H�/fi�q)�����y/�����͋ /�T���&0�&5 ��  ~e�j-�i;�芽����y&w&������ 4��&��Á����� ����FH?�q�6�/����6��6���??��y�&����4�ŀ�3�G�ݨ�����̀�%�.2����ˁ P    z	�n���щ,qqs��������g��,���;�t��lw/r(�!��5y�ό~�0�jt�{�~ fz��q��ek��ό ~B~�5i��~q& �/���c���D�6q!>&(?�/�7�/�:���wg)6 �{�:�/7�j:!.��/{�?��F�d��9F�J�)��)�-&.�f-(?�/�`��/�d�v�����l ?�B��/b������-�B. O�m�Țx)p���d0
  F������ �� �� �zi�-"(7���g��,����ڀ�q7�t��(������!/�eI��D� ����t&� �P�&/F.��F�, �7  ���0&� �k��� ��� ��/�˲l�t�	� ��à�����-�  `m�mޛ ��)����(� ���c�
F��4
c!�����J��K t	�f;-&.7f89fP0&
/f�h�x��
6�@.�/���P����
�"��
H.0�&
6B�����7��x6&��B���2@��Шa6�H?独�Ш7�J7-&8�* ��6��л ����	�J:0d��*CF�;T�`k�Ѝ��ch��q�����m�����ܨ/틬���z��# ���                                                                                                                                                                                                