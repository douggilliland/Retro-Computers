
--
-- Copyright (c) 2008-2019 Sytse van Slooten
--
-- Permission is hereby granted to any person obtaining a copy of these VHDL source files and
-- other language source files and associated documentation files ("the materials") to use
-- these materials solely for personal, non-commercial purposes.
-- You are also granted permission to make changes to the materials, on the condition that this
-- copyright notice is retained unchanged.
--
-- The materials are distributed in the hope that they will be useful, but WITHOUT ANY WARRANTY;
-- without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
--

-- $Revision: 1.16 $

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity vga is
   port(
      base_addr : in std_logic_vector(17 downto 0);

      bus_addr_match : out std_logic;
      bus_addr : in std_logic_vector(17 downto 0);
      bus_dati : out std_logic_vector(15 downto 0);
      bus_dato : in std_logic_vector(15 downto 0);
      bus_control_dati : in std_logic;
      bus_control_dato : in std_logic;
      bus_control_datob : in std_logic;

      vga_cursor : in std_logic_vector(12 downto 0);

      vga_hsync : out std_logic;
      vga_vsync : out std_logic;
      vga_out : out std_logic;

      reset : in std_logic;
      clk : in std_logic;
      clk50mhz : in std_logic
   );
end vga;

architecture implementation of vga is

signal base_addr_match : std_logic;

subtype u is std_logic_vector(7 downto 0);
type mem_type is array(0 to 2047) of u;

signal meme : mem_type;
signal memo : mem_type;

signal vgaclk : std_logic := '0';
signal vga_col : integer range 0 to 1039 := 0;
signal vga_row : integer range 0 to 665 := 0;
signal vga_fontcolumnindex : std_logic_vector(2 downto 0) := "000";
signal vga_fontrowindex : std_logic_vector(3 downto 0) := "0000";
signal vga_charindex : std_logic_vector(12 downto 0) := "0000000000000";
signal vga_rowstartindex : std_logic_vector(12 downto 0) := "0000000000000";

signal cursor_match : std_logic_vector(2 downto 0) := "000";
signal char_evn, char_odd : std_logic_vector(7 downto 0);
signal ix : std_logic_vector(14 downto 0);
signal fb : std_logic;
signal even_odd : std_logic;

constant vga_font : std_logic_vector(0 to 24575) :=
   "0001110111111000111111010101101100000000000000000000000000000000"  &   -- 0
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 64
   "0000000000000000000000000000000000000000000000010000000000000000"  &   -- 128
   "0000000000000000000000000000000000000000000000000000000001000000"  &   -- 192
   "1111111110001111111110111111111000000000000000000000000000000000"  &   -- 256
   "0000000000000000000000000000000000000000000000000000000000000001"  &   -- 320
   "0001101000010001010001100000100000000011010000110000100000000010"  &   -- 384
   "0000000000000000010101010101010110000000000010001010000001000000"  &   -- 448
   "1111111110001111111110111111111000000000000000000000000000000000"  &   -- 512
   "0000000000000000000000000000000000000000000000000000000000000001"  &   -- 576
   "1011111000110011011011100101100000000011011000110000100000100010"  &   -- 640
   "0000000000000000010101010101010110100100100010001010000000010000"  &   -- 704
   "1111111110001111111110111101111000000001000000000000000000000000"  &   -- 768
   "0000000000000000000000000000000010000000000000000000000000000000"  &   -- 832
   "1111011011101110011111000111000000000001011000110000000000100000"  &   -- 896
   "0101010101010101000000000000000001100100101000101000100000010000"  &   -- 960
   "1110000001011111000001111101100100000001000000000000000000000000"  &   -- 1024
   "0000000000000000000000000000000010000000000000000000000000000000"  &   -- 1088
   "0110111011111110000110100011110000000011011000110000100000100000"  &   -- 1152
   "0101010101010101010101010101010101000100010001101001000000100100"  &   -- 1216
   "1000000000000000000000000000000000000001000000000000000000000000"  &   -- 1280
   "0000000000000000000000000000000010000000000000000000000000000001"  &   -- 1344
   "0001101000010011010001100000110000000011011000110000100000000010"  &   -- 1408
   "0000000000000000010101010101010100000000010001000001000000100100"  &   -- 1472
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 1536
   "0000000000000000000000000000000000000000000000000000000000000001"  &   -- 1600
   "0001001000000001010001000000000000000000010000110000000000000010"  &   -- 1664
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 1728
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 1792
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 1856
   "0000000000000000000000000000000000000000000000010000000000000000"  &   -- 1920
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 1984
   "1111111111111111111111111111111100000000000000000000010100000000"  &   -- 2048
   "0010111010011110101001111010000000100000100110000000000000000000"  &   -- 2112
   "0001001000000000110001000000001000000001010000100000000000000000"  &   -- 2176
   "0000000000000000000000000000000000000000000000000000000000001011"  &   -- 2240
   "1000000000000000000001000000000000000000000000001011011111000011"  &   -- 2304
   "1010111110111111111111111111010000100000100110000000000000000111"  &   -- 2368
   "0011111000110011110011101001101100000101101000000000001010101010"  &   -- 2432
   "0000000000000000010101010101010100111100000100010100011001011011"  &   -- 2496
   "0000000000000000000000000010000000100010010000001011011111000011"  &   -- 2560
   "1111111101101001111110000111010000100000100110000000100000000111"  &   -- 2624
   "0110110101110111100110101011101100011110101000001011101011101010"  &   -- 2688
   "0000000000000000010101010101010111111100001110111110111001010010"  &   -- 2752
   "0000000000000000000000000000000001101011010000001111011111000001"  &   -- 2816
   "1111111101101001111110000011011010001010010010000000100000001110"  &   -- 2880
   "1101001101000100111101001110011100011010000000001011101001000000"  &   -- 2944
   "0101010101010101000000000000000011110000111011101111110000110110"  &   -- 3008
   "0000001111010000111111000000001101000011100000001111111111001001"  &   -- 3072
   "1111111101100001111110000011011010001010011000000000000000011000"  &   -- 3136
   "1011111110111000111011101101110100011010101000001011101010101000"  &   -- 3200
   "0101010101010101010101010101010100101100111101110001101000111100"  &   -- 3264
   "0000000000000000000000000000000000100001100000001011111111001001"  &   -- 3328
   "1011011111010111111111111111010010001010001000000000000000010011"  &   -- 3392
   "0011110110111011010011101001100100001101101000000000001010101010"  &   -- 3456
   "0000000000000000010101010101010100011100000100110100011000001001"  &   -- 3520
   "1000000000000000000000000000000000100000000000000000010100000000"  &   -- 3584
   "0000011010010110000011111110000000000000000000000000000000010011"  &   -- 3648
   "0000000000000011000000001000000000000101000000000000001000001010"  &   -- 3712
   "0000000000000000000000000000000000010000000000000100010000000001"  &   -- 3776
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 3840
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 3904
   "0000000000000000000000000000000000000000010000100000001000000000"  &   -- 3968
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 4032
   "1001111111101100111111011101111100000000000000001011011111000001"  &   -- 4096
   "1000000110010111010101111010000000000000000000000000000000000010"  &   -- 4160
   "0000001000000000000000001000000100000001010000100000001000001000"  &   -- 4224
   "1000000000000000000000000000000000110000000000000100010000011001"  &   -- 4288
   "0111111111011011000000110101101000001010000000001111011111000001"  &   -- 4352
   "1111111110011111111111111111000000100000100100000000000000000010"  &   -- 4416
   "0000001100000000100000001000001100011101001000001011001001101000"  &   -- 4480
   "1000000000000000010101010101010101111000001100111100111000011011"  &   -- 4544
   "0111111111001011000001110111101000101010000000000100000000000010"  &   -- 4608
   "0111111000001010101000000101001000100010100110000000100000000000"  &   -- 4672
   "0010010100000000100000000000001000011100101000101011000011100000"  &   -- 4736
   "1000000000000000010101010101010101001100011101111001101001100110"  &   -- 4800
   "1110001111010011000000100000111001101000110000000100100000001010"  &   -- 4864
   "0000000001100000000010000000001010000010010010000000100000011110"  &   -- 4928
   "0010011000000000000000000000000000100000110000100000001011001000"  &   -- 4992
   "1101010101010101000000000000000010010100010011001111010101100100"  &   -- 5056
   "1000001001000000111111000000010101001011110000000100100000001000"  &   -- 5120
   "0100100001110000000010000000011010001000011000000000000000011110"  &   -- 5184
   "0010011000000000100000000000000000010000111000101011001010101000"  &   -- 5248
   "1101010101010101010101010101010110111100101110011110111100011000"  &   -- 5312
   "0000000000000000000000000000000000101011000000001011101111000001"  &   -- 5376
   "1111111110010111111101111110011000001010001000000000000000000010"  &   -- 5440
   "0000000100000000100000001000000100010101001000001011000000100000"  &   -- 5504
   "1000000000000000010101010101010100111000101100110100111000011001"  &   -- 5568
   "0000000000000000000000000000000000100000000000001011001111000001"  &   -- 5632
   "1011011110000111111111111110000000000010000000000000000000000000"  &   -- 5696
   "0000000100000000000000001000000100001101000000000000001000001000"  &   -- 5760
   "1000000000000000000000000000000000000000000000100000000000000001"  &   -- 5824
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 5888
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 5952
   "0000000000000000000000000000000000000000010000100000001000001000"  &   -- 6016
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 6080
   "1001111111101100111111011101111100001000000000001010011011000001"  &   -- 6144
   "1101000110010111010101110010100000000000000000000000000000000000"  &   -- 6208
   "0000001111110000010000001111100100000000010000100000101000011000"  &   -- 6272
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 6336
   "0000000000010000000000000000000000011100001000001010011011000001"  &   -- 6400
   "1111111110011111111101111101101000100000100100000000000000000001"  &   -- 6464
   "0000001111110000111111101111111100111011000000000000101000011010"  &   -- 6528
   "0000000000000000010101010101010100000011000000000000000000000010"  &   -- 6592
   "0000000000000000000000000010001000010110101000000000100000001000"  &   -- 6656
   "0010111000001110101000001101001000100010100110000000100000000001"  &   -- 6720
   "1101100011111111101111100000011000111111011100101000100001100011"  &   -- 6784
   "0000000000000000010101010101010100000011000000000000000000000010"  &   -- 6848
   "1000000000010000000001000000000001101011100100000100100000001010"  &   -- 6912
   "0000000001110000000010000000000000000010000010000000100000011100"  &   -- 6976
   "1101101011111111001111100000001001100110001100001111101001111001"  &   -- 7040
   "0101010101010101000000000000000000000011000000000000000100000000"  &   -- 7104
   "1110001111000011111111100000010101010011011100000100100100110010"  &   -- 7168
   "0000000001110100000010001010010010001000000000000000000000011100"  &   -- 7232
   "1101101011111111001111101000001001100110001000001111101000111000"  &   -- 7296
   "0101010101010101010101010101010100000011000000001000000100000000"  &   -- 7360
   "0000000000000000000000000000000000111000011000011011100111110001"  &   -- 7424
   "1110100110000111111001111110011010001000000000000000000000000001"  &   -- 7488
   "0000000011111111111111101111111100100110011100100000100000000010"  &   -- 7552
   "0000000000000000010101010101010100000011000000001000000000000000"  &   -- 7616
   "0000000000000000000000000000000000001100000000011011000011000001"  &   -- 7680
   "1110100110000111111001110100001000000000000000000000000000000001"  &   -- 7744
   "0000000011110000110000001111110100000000001100000000101000001010"  &   -- 7808
   "0000000000000000000000000000000000000010000000000000000000000000"  &   -- 7872
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 7936
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 8000
   "0000000000000000000000000000000000000000010000100000001000001000"  &   -- 8064
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 8128
   "1111111111101011111111110111101000010000000000001000011011000100"  &   -- 8192
   "1101000110010111010001110000000000000000000000101010111111100000"  &   -- 8256
   "0000001100000000011111101111100100101010010000100000111010001000"  &   -- 8320
   "0000000000000000000000001111111100000011000000000100000001111101"  &   -- 8384
   "1111110110100111111110111111010100011100000000001000111011001100"  &   -- 8448
   "1111111110011111111101110101100001111101110101111111111111100001"  &   -- 8512
   "1111111111110000111111111111111100111011100100000001111010011110"  &   -- 8576
   "0000000000000000010111111111111111111111111100001111111011111111"  &   -- 8640
   "1111110110110111111110111111010100011110101000000000100000001100"  &   -- 8704
   "0010111000011110101100001101100001111111110111010101100000100001"  &   -- 8768
   "1111110011110000110000010000011000011001110100100011000011010111"  &   -- 8832
   "0000000000000000011111111111111111111100111111111011111010000010"  &   -- 8896
   "1111110110100111111110111111011101011010101100000100000100000100"  &   -- 8960
   "1000000001110110000010001010000001111111011010111111100000111100"  &   -- 9024
   "0010011000001111000000001000000001101101100000000110001011001001"  &   -- 9088
   "0101010101010101001010101010101011111110111111111111111010000010"  &   -- 9152
   "0000001001100100000001011111000001010010011100010110100100110111"  &   -- 9216
   "1000000001100100000010001010010001111100111001111011110000111100"  &   -- 9280
   "1111111000001111000000011000000001001101100100000101011010011100"  &   -- 9344
   "0101010101010101011111111111111111111110111111111111111011111010"  &   -- 9408
   "0000000000000000000000000000000000010100010000011011100011110111"  &   -- 9472
   "1110100010000111111001110100010000111101101101111111111111100001"  &   -- 9536
   "1111110011110000111111111111111100100011100100100001110010011110"  &   -- 9600
   "0000000000000000011111111111111100000001111100001111111011111101"  &   -- 9664
   "1000000000000000000000000000000000010100000000001001000011000100"  &   -- 9728
   "1110100010000111111001110100000000000001000100000100001111100001"  &   -- 9792
   "0000000011110000111111101111111100100010000000000000101010001010"  &   -- 9856
   "0000000000000000001100110011001100000011000000001000000010000101"  &   -- 9920
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 9984
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 10048
   "0000000000000000000000000000000000000000010000100000001000001000"  &   -- 10112
   "0000000000000000001100110011001100000010000000000000000000000000"  &   -- 10176
   "1000000000000000000000000000000000000000001001001000111000001000"  &   -- 10240
   "1101000110010111010001110000000000011111000001010101011101100000"  &   -- 10304
   "1111111100000000111111101111100100110011110100100000010010001100"  &   -- 10368
   "0000000011111111000000000000000000000001111100001011111011111101"  &   -- 10432
   "1000000000000000000000000000000000010010001101001000111011001000"  &   -- 10496
   "1111111110011111111001110001000000111111100101111111011111010001"  &   -- 10560
   "1111111111110000111111101111111100111111101111000110011001101100"  &   -- 10624
   "0000000011111111010111110000000000000001111100001111111111111111"  &   -- 10688
   "1000000000000000000000000000000000011010101101000001011111000000"  &   -- 10752
   "0010111010011000101100001111100000100010100111101010100010010001"  &   -- 10816
   "0000001011110000110000010000011000011100011011100111001001110010"  &   -- 10880
   "0000000011111111011111110000000000000000000000000100000100000010"  &   -- 10944
   "0000000000000000000000000000000001001010101101011111011111000001"  &   -- 11008
   "1010011011110110101110011110100000000010110011000000100000011000"  &   -- 11072
   "0000001000001111110000011000000000110100001111100111001101111110"  &   -- 11136
   "0111111111111111001000000000000000000010000011110000000100000000"  &   -- 11200
   "0000000000000000000000000000000001011100011101010111111011000001"  &   -- 11264
   "1010011011100000101110001100010001001011011101000100010010101100"  &   -- 11328
   "0000001000001111000000010000000100000100001111100111111111101110"  &   -- 11392
   "0111111111111111010011001100110011111110000011110000000111111010"  &   -- 11456
   "1000000000000000000000000000000000010100011101001001111011000010"  &   -- 11520
   "1110111010000111111001110100010001111111101101111111011111100101"  &   -- 11584
   "1111111000000000111111101111111100000101101011000110110010110010"  &   -- 11648
   "0011001100110011010011001100110011111100111100001111111111111111"  &   -- 11712
   "1000000000000000000000000000000000000010001101001000000001000010"  &   -- 11776
   "1100100010000111010001110000000000110101100001111011001101000101"  &   -- 11840
   "1111111000000000111111101111111000000101101011000100001000010100"  &   -- 11904
   "0011001100110011000000000000000000000010111100001111111110000101"  &   -- 11968
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 12032
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 12096
   "0000000000000000000000000000000000000000010000100000001000000000"  &   -- 12160
   "0011001100110011000000000000000000000010000000000000000000000000"  &   -- 12224
   "1000000000000000000000000000000000000010000000001000101010000100"  &   -- 12288
   "1101000110010111010001110000000000011101000001010100011101000000"  &   -- 12352
   "1111111100000000011111101111100100101001010000100000010000001100"  &   -- 12416
   "0000000000000000000000001111111100000001111100001011111011111101"  &   -- 12480
   "1000000000000000000000000000000000010010000000001000101010001100"  &   -- 12544
   "1111111110011111111001110011000001111101100101111111011101000000"  &   -- 12608
   "1111111111110000111111101111101100111011100100000000010000011100"  &   -- 12672
   "0000000000000000010111111111111111111111111100001111111011111111"  &   -- 12736
   "1000000000000000000000000000000000010010101000010010100100001100"  &   -- 12800
   "0110111000001000101000011011000001100110100110101011100010000001"  &   -- 12864
   "0000000011110000100000011000011000011010110100100000100000010001"  &   -- 12928
   "0000000000000000011111111111111111111110111100000100000000000010"  &   -- 12992
   "0111100001111100000100111100000001001110101100010110100100000101"  &   -- 13056
   "1100000001110010001010011100100001000110010111000001100110111101"  &   -- 13120
   "0000001011111111010000011000010001101110100000000100101110001111"  &   -- 13184
   "0000111100001111011100001111000011111110111111110000000010000000"  &   -- 13248
   "0000111111111111111101010010111101011110011100000100100000000111"  &   -- 13312
   "1100000101110010001110011100110001001100011100000100010010111101"  &   -- 13376
   "0000001011111111010000010000010001001110000100000100111110011110"  &   -- 13440
   "0000111100001111011111111111111111111110111111110000000011111010"  &   -- 13504
   "1000110011111111011110010011111100011010010000001001111011000110"  &   -- 13568
   "1110100110000111010101110000010001101101101001111100011101000001"  &   -- 13632
   "1111110111110000111111101111111100000011010110100000010000010100"  &   -- 13696
   "0000000000000000011111111111111111111110111100001111111011111111"  &   -- 13760
   "1000110011111111000010010011111100000010000000001001111011000100"  &   -- 13824
   "1110100110000111010001110000000000100101100001111000001101000000"  &   -- 13888
   "1111110100000000111111101111101100000001000010000000001000000100"  &   -- 13952
   "0000000000000000001100110011001100000010111100001111111010000101"  &   -- 14016
   "1111101011111000000001101101111100000000000000000000000000000000"  &   -- 14080
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 14144
   "0000000000000000000000000000000000000000010000100000001000000000"  &   -- 14208
   "0000000000000000001100110011001100000010000000000000000000000000"  &   -- 14272
   "1000000000000000000000000000000000001010000000001000001010000000"  &   -- 14336
   "1101000110110111010001010010000001011101000001010100010101000000"  &   -- 14400
   "1111111000000000011111101111100100100000010000100000010000011100"  &   -- 14464
   "0000000000000000100000000000000011111111111100001011111011111101"  &   -- 14528
   "1000000000000000000000000000000000011010001000011010001010000000"  &   -- 14592
   "1111111110011111111001111011000001111101100101111110011101000000"  &   -- 14656
   "1111111111110000111111111111101100111001000000000000110000011100"  &   -- 14720
   "0000000000000000100011110000111111111111111100001111111011111111"  &   -- 14784
   "1000000000000000000000000000000000010100101000010010000100001000"  &   -- 14848
   "0010111000001000101000111001000000100010100110101010101010100000"  &   -- 14912
   "1111110111110000100000011000001000011101000100100000100010000001"  &   -- 14976
   "0000000000000000100011110000111100000000000000000100000010000010"  &   -- 15040
   "1100010010101110011000011110111101001100100100000100000100001010"  &   -- 15104
   "1000000001100000000010000100000000000010010011000001100110111101"  &   -- 15168
   "1111111000001111000000000000011001100101110100000100001010011111"  &   -- 15232
   "0000111100001111100000000000000000000010000011110000000110000000"  &   -- 15296
   "1011001100000000100011101101000001010010011110000100100000110010"  &   -- 15360
   "1000000001110010001010111100110001001000011100000101011011011101"  &   -- 15424
   "1111111000001111010000010000011001000101110000000100011000011110"  &   -- 15488
   "0000111100001111100011110000111111111110000011110000000101111111"  &   -- 15552
   "1000100001010001010000000000000000011010011010001001111011110000"  &   -- 15616
   "1110100110010111011101111000110001101001101101111101011101000000"  &   -- 15680
   "1111110100000000111111111111101100110111100110100000010000000000"  &   -- 15744
   "0000000000000000100011110000111111111101000000001111111011111111"  &   -- 15808
   "1011001000000000001111100100000000001000000000001001011011000000"  &   -- 15872
   "0110100110001111010101010010000000100001100001111000000101000000"  &   -- 15936
   "1111110100000000111111101111100100110010000110000000101000000000"  &   -- 16000
   "0000000000000000100000000000000000000001000000001111111010000101"  &   -- 16064
   "1100010000000110000000011110000000000000000000000000000000000000"  &   -- 16128
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 16192
   "0000000000000000000000000000000000000000010000100000001000001000"  &   -- 16256
   "0000000000000000100000000000000000000000000000000000000000000000"  &   -- 16320
   "1000000000000000000000000000000000010010000000011011011011000000"  &   -- 16384
   "1100000110110111010101011010000001011100000001010001010100000000"  &   -- 16448
   "1111111000000000011111101111100100010010110000100000110000001100"  &   -- 16512
   "0000000000000000000000000000000011111110111100001011111011111000"  &   -- 16576
   "1000000000000000000000000000000000011110000000011011011011000000"  &   -- 16640
   "1111111110111111111101011011000001111101100101111111010111100000"  &   -- 16704
   "1111111011110000111111101111101100111010100000000000110010001101"  &   -- 16768
   "0000000000000000000011110000111111111111111100001111111011111111"  &   -- 16832
   "1000000000000000000000000000000000011100000000000000000100000010"  &   -- 16896
   "0011111000001000101000100001000000100011100110101110101111100000"  &   -- 16960
   "0000000111110000100000000000001001111000000000000000000010000001"  &   -- 17024
   "0000000000000000000011110000111100000001000000000100000010000111"  &   -- 17088
   "0100010000101110000010011110000000011000110000100100000100001011"  &   -- 17152
   "0000000001100000010010100100000001000011010010001100101101011101"  &   -- 17216
   "0000001100001111000000000000010101110100000000000000001000001110"  &   -- 17280
   "0000111100001111000000000000000011111111000011110000000100000111"  &   -- 17344
   "0100001110101100100011010011111100011010110010100100100000111001"  &   -- 17408
   "0000100001100010000010100100010001001001011000001100011110011101"  &   -- 17472
   "0000001100001111100000000000010001100101000000000000011000001110"  &   -- 17536
   "0000111100001111000011110000111111111111000011110000000101111010"  &   -- 17600
   "1111101011111101011111111110111100011110000010001011111011110000"  &   -- 17664
   "0111110110011111011101011010110001111101101101111101010111000000"  &   -- 17728
   "1111110111110000111111101111100101110011100010000000110000001000"  &   -- 17792
   "0000000000000000000011110000111111111101111100001111111011111101"  &   -- 17856
   "1100000010000100000010010010111100010100000000001011011011000000"  &   -- 17920
   "0111010110011111011101011010100000110101100101110001000101100000"  &   -- 17984
   "1111110011110000011111101111100100011010100010000000101010001100"  &   -- 18048
   "0000000000000000000000000000000000000010111100001111111010000101"  &   -- 18112
   "1100010000000110000000001110000000000000000000000000000000000000"  &   -- 18176
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 18240
   "0000000000000000000000000000000000000000010000100000001000001000"  &   -- 18304
   "0000000000000000000000000000000000000010000000000000000000000000"  &   -- 18368
   "1000000000000000000000000000000000000100000000000010000000000000"  &   -- 18432
   "0110111010011110101000011010000000100000101111000010000010100000"  &   -- 18496
   "1111111011110000110000001000001110000001000000000000110010000001"  &   -- 18560
   "0000000000000000000000000000000000000000000000000000000010000000"  &   -- 18624
   "1000000000000000000000000000000000010110000000001111011011000010"  &   -- 18688
   "1110111110111111111101011011010001111110111111111011010110100100"  &   -- 18752
   "1111111011110000111111101111101100010011110000100100110010001101"  &   -- 18816
   "0000000000000000000011110000111111111110111100001111111011111010"  &   -- 18880
   "1000000000000000000000000000000000010010010000001111011111000010"  &   -- 18944
   "1011111101101001111111000111010001111110110110111011010100100101"  &   -- 19008
   "0000000011111111101111101111111001011010110000100100110010001110"  &   -- 19072
   "0000000000000000000011110000111111111110111111111111111011111010"  &   -- 19136
   "0100010000101110000000011110000001001010010000101111011111000001"  &   -- 19200
   "1011111101101001110111100111010001111110010010010011111000101101"  &   -- 19264
   "0000001111111111101111101111111101101110110000100100111010000010"  &   -- 19328
   "0000111100001111000000000000000011111111111111111011111011111000"  &   -- 19392
   "0011001100000000101001000001000001010000100010101111111011011001"  &   -- 19456
   "1011110101001001010111000111010000111110011010010101100100111001"  &   -- 19520
   "0000001111111111101111101111110101011110110000100100101010001110"  &   -- 19584
   "0000111100001111000011110000111100000011111111111011111010000000"  &   -- 19648
   "1000100001010001010000100000000000010110100010001111111011011000"  &   -- 19712
   "1111010111011111011111011111010001111101111111110101110111110001"  &   -- 19776
   "1111111011111111011111101111110101011011110000100100110010001111"  &   -- 19840
   "0000000000000000000011110000111111111110111111111111111011111101"  &   -- 19904
   "1011011000000100000111001000000000000110000000000110000000000000"  &   -- 19968
   "1100010010011110001000011010000001001001110101100000010011110000"  &   -- 20032
   "1111111011110000010000000000000010000001010000100100111010001001"  &   -- 20096
   "0000000000000000000000000000000011111110000000000100000001111101"  &   -- 20160
   "1100010010000010000000011110111100000000000000000000000000000000"  &   -- 20224
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 20288
   "0000000000000000000000000000000000000000000000000000001000000000"  &   -- 20352
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 20416
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 20480
   "0000000000000000000000000000000000000001001000000000000001000000"  &   -- 20544
   "0000000100000000000000000000000110000001000000000000010000000001"  &   -- 20608
   "0000000000000000000000000000000000000000000000000000000000000101"  &   -- 20672
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 20736
   "0000000000000000000000000000000000000001001000001000000001000000"  &   -- 20800
   "0000000100000000000000000000000010000001000000000000010000000001"  &   -- 20864
   "0000000000000000000011110000111100000001000000000000000000000111"  &   -- 20928
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 20992
   "0000000000000000000000000000000000000000000000001000000000000000"  &   -- 21056
   "0000000000000000000000000000000011000000000000000000000000000000"  &   -- 21120
   "0000000000000000000011110000111100000001000000000000000000000010"  &   -- 21184
   "1111000010101100011100011110111101000000000010000000000000010000"  &   -- 21248
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 21312
   "0000000000000000000000000000000011000000000000000000000000000000"  &   -- 21376
   "0000111100001111000000000000000000000000000000000000000000000000"  &   -- 21440
   "1000011110000011111101010000111101000000000010000000000000010000"  &   -- 21504
   "0000000000000000000000000000000000000000001000000100000000000000"  &   -- 21568
   "0000000100000000000000000000000011000000000000000000000000000000"  &   -- 21632
   "0000111100001111000011110000111100000001000000000000000000000000"  &   -- 21696
   "1000110111010011111100110001111100000000000000000000000000000000"  &   -- 21760
   "0000000000000000010000000000000000000001001000000100000001000000"  &   -- 21824
   "0000000100000000000000000000000011000001000000000000000000000001"  &   -- 21888
   "0000000000000000000011110000111100000001000000000000000000000101"  &   -- 21952
   "1000010110000011111010010001111100000000000000000000000000000000"  &   -- 22016
   "0000000000000000010000000000000000000001000000000000000001000000"  &   -- 22080
   "0000000000000000000000000000000010000001000000000000000000000001"  &   -- 22144
   "0000000000000000000000000000000000000000000000000000000000000101"  &   -- 22208
   "0111001100000100110001001111000000000000000000000000000000000000"  &   -- 22272
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 22336
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 22400
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 22464
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 22528
   "0000000000000000000000000000000100000000000000001000000000000000"  &   -- 22592
   "0000000000000000000000000000000000000000000000000000010000000000"  &   -- 22656
   "0000000000000000000000000000000000000000000000000000000000000010"  &   -- 22720
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 22784
   "0000000000000000000000000000000100000001001000001000000001000000"  &   -- 22848
   "0000000000000000000000000000000000000001000000000000010000000001"  &   -- 22912
   "0000000000000000000011110000111100000000000000000000000000000111"  &   -- 22976
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 23040
   "0000000000000000000000000000000100000001001000001000000001000000"  &   -- 23104
   "0000000100000000000000000000000000000001000000000000000000000001"  &   -- 23168
   "0000000000000000000011110000111100000001000000000000000000000111"  &   -- 23232
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 23296
   "0000000000000000000000000000000100000001001000001100000001000000"  &   -- 23360
   "0000000100000000000000000000000001000001000000000000000000000001"  &   -- 23424
   "0000111100001111000000000000000000000001000000000000000000000111"  &   -- 23488
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 23552
   "0000000000000000000000000000000100000001001000000100000001000000"  &   -- 23616
   "0000000100000000000000000000000001000001000000000000000000000001"  &   -- 23680
   "0000111100001111000011110000111100000001000000000000000000000101"  &   -- 23744
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 23808
   "0000000000000000000000000000000100000001000000000100000001000000"  &   -- 23872
   "0000000000000000000000000000000000000001000000000000000000000001"  &   -- 23936
   "0000000000000000000011110000111100000000000000000000000000000101"  &   -- 24000
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 24064
   "0000000000000000000000000000000100000000000000000100000000000000"  &   -- 24128
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 24192
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 24256
   "0000010000000000000000000000000000000000000000000000000000000000"  &   -- 24320
   "0000000000000000000000000000000100000000000000000000000000000000"  &   -- 24384
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 24448
   "0000000000000000000000000000000000000000000000000000000000000000"   -- 24512
;


begin
   base_addr_match <= '1' when base_addr(17 downto 13) = bus_addr(17 downto 13) else '0';
   bus_addr_match <= base_addr_match;

   process(clk50mhz)
   begin
      if clk50mhz = '1' and clk50mhz'event then
         if reset = '1' then
            vgaclk <= '0';
         else
            vgaclk <= not vgaclk;
         end if;
      end if;
   end process;

   process(clk, base_addr_match)
   begin
      if clk = '1' and clk'event then
         bus_dati(7 downto 0) <= meme(conv_integer(bus_addr(12 downto 1)));
         bus_dati(15 downto 8) <= memo(conv_integer(bus_addr(12 downto 1)));

         if base_addr_match = '1' and bus_control_dato = '1' then
            if bus_control_datob = '0' or (bus_control_datob = '1' and bus_addr(0) = '0') then
               meme(conv_integer(bus_addr(12 downto 1))) <= bus_dato(7 downto 0);
            end if;
            if bus_control_datob = '0' or (bus_control_datob = '1' and bus_addr(0) = '1') then
               memo(conv_integer(bus_addr(12 downto 1))) <= bus_dato(15 downto 8);
            end if;
         end if;
      end if;
   end process;

   process(vgaclk)
   begin
      if vgaclk='1' and vgaclk'event then
         if reset = '1' then
            vga_col <= 0;
            vga_row <= 0;
            vga_rowstartindex <= "0000000000000";
            vga_fontrowindex <= "0000";
            vga_hsync <= '1';
            vga_vsync <= '1';
            vga_out <= '0';
         else
            if vga_col < 799 then
               vga_col <= vga_col + 1;
            else
               vga_col <= 0;
               if unsigned(vga_fontrowindex) < unsigned'("1011") then
                  vga_fontrowindex <= vga_fontrowindex + 1;
               else
                  vga_fontrowindex <= "0000";
                  vga_rowstartindex <= vga_rowstartindex + 80;
               end if;
               if vga_row < 523 then
                  vga_row <= vga_row + 1;
                  if vga_row >= 479 then
                     vga_rowstartindex <= "0000000000000";
                     vga_fontrowindex <= "0000";
                  end if;
               else
                  vga_row <= 0;
                  vga_rowstartindex <= "0000000000000";
                  vga_fontrowindex <= "0000";
               end if;
            end if;

            vga_hsync <= '1';
            vga_out <= '0';

            if (vga_charindex = vga_cursor) then
               cursor_match <= cursor_match(1 downto 0) & '1';
            else
               cursor_match <= cursor_match(1 downto 0) & '0';
            end if;

            if vga_charindex(0) = '0' then
               even_odd <= '0';
            else
               even_odd <= '1';
            end if;
            char_evn <= meme(conv_integer(vga_charindex(12 downto 1)));
            char_odd <= memo(conv_integer(vga_charindex(12 downto 1)));
            if even_odd = '0' then
               ix <= (vga_fontrowindex & "00000000000") + (vga_fontcolumnindex & "00000000") + char_evn;
            else
               ix <= (vga_fontrowindex & "00000000000") + (vga_fontcolumnindex & "00000000") + char_odd;
            end if;
            fb <= vga_font(conv_integer(ix));

            if vga_col < 96 then
               vga_hsync <= '0';
            elsif vga_col < 141 then
               vga_fontcolumnindex <= "111";
               vga_charindex <= vga_rowstartindex;
            elsif vga_col < 784 then

               if unsigned(vga_fontcolumnindex) = unsigned'("110") then
                  vga_charindex <= vga_charindex + 1;
               end if;

               if unsigned(vga_fontcolumnindex) < unsigned'("111") then
                  vga_fontcolumnindex <= vga_fontcolumnindex + 1;
               else
                  vga_fontcolumnindex <= "000";
               end if;

               if vga_col < 144 then
                  vga_out <= '0';
               else
                  vga_out <= fb;
               end if;

               if cursor_match(2) = '1' then
                  vga_out <= '1';
               end if;

            end if;

            vga_vsync <= '1';
            if vga_row < 480 then                                              -- 480 normal display rows
            elsif vga_row < 489 then                                           -- 10 rows - front porch
               vga_out <= '0';
            elsif vga_row < 491 then                                           -- 2 rows - sync pulse
               vga_vsync <= '0';
               vga_out <= '0';
            else                                                               -- 33 rows - back porch
               vga_out <= '0';
            end if;

         end if;
      end if;
   end process;

end implementation;

