���    �# :		4(*;:  8 8 2 > 
-	" :6"
5.* 0 2	%9
032?
    
>.
? 8   ( / :
+	)%!($  :       
 	* ( 4 2 +/47? % . % 	3
  8 
                                                                                                                                                                                                                                                                         ;` H	  h
�v
                                    `
            &    
  	  H	c	                                XR`MgSig�&�+�	1	�:  s1�	��u�	�'	,	�? ��A� ���   � @ � �����8	 �   ? �	���O	�""��H	�V	A\	E	�BE	����M	L	I	�	���
  ��
�\	)P	�M	����
.�-�
�O	�Z	_	����E	  R	���
H�J�;b	K	M	H�
�
D	_	~ �
�
!�J���
)(X	\	HM	@)���}M	�: 
�* $% �`
  F�(D������F��(�  D���| ���| J
�

��  | ��{ ���  �����z �(�. �!�
�E	A�
N!H�Fy	!%��
��D	���  �"""�  """��H	�  �A�C	��
  @@p���D	����C	����
�C	���%��
[	![	$S	$�F[	a@p���
$!%��
�$�
�$$�
��
  ${ x�����
  [	@�
��E	��H�
(FP%''��H	%&'%�&!$��
 && ''&{ �'| �'�
�	�$�(F!a$�S	&$'�%!&��
&{ �'| �'&'�
'%�
� �`   [	!�T	�w�Y	�
I	Z���
H	���$��
��h�
!�${ ���
$��% $��
$����
 �
���$�
�
@�
�
K	�
�${ `	 �
�BF�F�B�B�
U	��
�!$4�$E	:BE	�v�v���!%��
��
�y	�
      �
�  �u�
���F�D�@�!�������
E	n%�
�G	���
�G	���
$�
��}�t����F� �
 � ��
!����
�
  ��]	  �
�J�A\	�V	\	��L	M	�
�K	�
V	�
V	[	<<<<�
�
)��
s�22�F    �u _	 � �	$ ��1
��O	F�
�tFE	��${ �� �
E	�!J�$�${ ��@-FE	��
  .M	-M	�  ������2�]	  �(�
��	X�4��
��	���Y	v  ��
  ���H�
q��
���H�
������_	~ �
 F  r@� q�� 0 ����
[	!�E	�%��
+N	 :P	��;a ��
E	��
F  E	����� ��!]	 V�	H	��
�z �  ��
FV	�\	��3�
  �
$E	�$$S	` ����
�H	��
Q	> c	�
�
�v(H	 v�0F  �G	  �� (�X	�M	��
$'�'`%�'{ ��%$� a%��
=�
@
@@z

��7	 �  ��
�
����=�� ��
���| | J
J
 z  �(�
�(�
�(�
+�3%| 3%3�%x���
�FH	 1
�F  K	I	 k��8 e ���  �R	���!�
�&��  I	* J�w ��
���q��  ��
st�-�
�} t�  ����
�  3W	(<'<a3�
(�
)((��H	)&()(&!'��
 &&�((&P	X	�
'()!'��
'P	X	'�
()3<#Z	W	�0  T	 !Y	��
E	A�	�  7 ��%	�^ �  (9!(�<�
<<<(�
(�  �;a ��
 :P	��  M	� �(�"�H	D	 D	D	D	Z	�
  ##W	(:<;�   �
_	99`	H	9rH}-9W	�C G N L A B E `	������1
_	I	J @	
�D�F��Q	' �Jc	vK	���J������$�� �	 �U	 Q	! ��:((P	!3Y	�
3��
(�
30��
c	v    ��b	�_	I	� �
K	�
K	�U	U	E	��
�
_	I	[	��
K	��
��
��H�	�
����    ! > < " ^ @  	   E F I N O  S _ Q U X G M % ��
����om�������������������Y�V	U	!  \	! b	Y	�
X	�
c	v  ��E	�~M	� ���
�	���  !��_	I	X	 	
�
�F�  U	4!:( a!334 �
E	��
(P	��(3�
v  �$| �$�$�    V	< 3<E	��
  �
R	z (�
I	�	�z �  z ��E	���� ;,��E	 ��'�'���'���p	     � '�8��	6�5��� �����N����
  p��
�	�	��>���
�6	 	�
  �
�
����?�>�
�HNH	���    �    �!�| !X��DF�P�0�!�!��        �  �j��k�t�^<��7�=����@<�v  ���
���� ���Y	�
I	I%`	H	�t��
�H�^	~ �
F����
� ��
���
(�
 �X ��
. : ���	�������p	   ��p	       �
�� ��
��p	      �
���  ���
HNE	�H	  %qM	 : &> z  >�3�N	3�
5���6��	8��
���5p	 �  �
�������}} ��6	�   �
5�p	 �  HN�p		 v  ^	@u@x@�@����  F| ???�  43�!@4�
43�
�3���v�
�@���$g>�
.	��T   �
�
t ���  M	�         ���$!E	��$$E	�$!'$$!'� ���
��z �(/�`�
(�
�(�
Ps(�
�
�������
���� a� �> ��
�
�
� } ��F�/� �
�
ED�� a�� ����� w �,)  �� >@   8 �?��	��v
V  8 �! @ (( @    �^	�A S	iR�?z
�F�#	(V
�R
��  �	   ���" -?�?	�
�^��	e?	$^�?��! b>?� � ?�?��?	$�� ?	fQ
�	 ? �~ ��3��c	i   F   � >�                                                                �
'a	F  ��  ��    �
K	�  ��
E	��
+N	E	R	��V	<1
<F  �%� Z���	 �X C F R W B G   @  ��d 
 >A� ���7?� � � � � � ���7K����     ?  V	�G	#     "!9Z	F  a%H	!%�} ~ �G	  ! F  �
��E	��
  K	^	�                                                                                                                                                & ��	I	 ;���;�4�	�	�	�		 �� 	 O	 � �	 	 	 ��	 	 �	 �	JX�	 �������k�������������L��	 �q� ���*I^�/����	l����Q�F		 �	��	 	 � k                    { �(�(�  ����{ ��
�
���  ���
��p�&�p���a �  ��
���� t��
����� ����
{�������
� ��X	��
����  ��
��  (����
ia	�a	
 	��   
  ij 
4�H���
��
��%�Q	s��� �  �� $��
  8 ��
�
�y�