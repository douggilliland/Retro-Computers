library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sdbootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end sdbootstrap_ROM;

architecture arch of sdbootstrap_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"7f",
     2 => x"00",
     3 => x"00",
     4 => x"00",
     5 => x"00",
     6 => x"00",
     7 => x"08",
     8 => x"4f",
     9 => x"f9",
    10 => x"00",
    11 => x"7f",
    12 => x"00",
    13 => x"00",
    14 => x"70",
    15 => x"00",
    16 => x"30",
    17 => x"39",
    18 => x"81",
    19 => x"00",
    20 => x"00",
    21 => x"2a",
    22 => x"c0",
    23 => x"fc",
    24 => x"03",
    25 => x"e8",
    26 => x"80",
    27 => x"fc",
    28 => x"04",
    29 => x"80",
    30 => x"33",
    31 => x"c0",
    32 => x"81",
    33 => x"00",
    34 => x"00",
    35 => x"02",
    36 => x"46",
    37 => x"fc",
    38 => x"27",
    39 => x"00",
    40 => x"33",
    41 => x"fc",
    42 => x"f0",
    43 => x"00",
    44 => x"81",
    45 => x"00",
    46 => x"00",
    47 => x"06",
    48 => x"33",
    49 => x"fc",
    50 => x"00",
    51 => x"01",
    52 => x"81",
    53 => x"00",
    54 => x"00",
    55 => x"04",
    56 => x"41",
    57 => x"fa",
    58 => x"00",
    59 => x"72",
    60 => x"61",
    61 => x"00",
    62 => x"02",
    63 => x"d6",
    64 => x"33",
    65 => x"fc",
    66 => x"0f",
    67 => x"00",
    68 => x"81",
    69 => x"00",
    70 => x"00",
    71 => x"06",
    72 => x"2e",
    73 => x"3c",
    74 => x"00",
    75 => x"00",
    76 => x"07",
    77 => x"ff",
    78 => x"41",
    79 => x"f9",
    80 => x"80",
    81 => x"00",
    82 => x"08",
    83 => x"00",
    84 => x"10",
    85 => x"fc",
    86 => x"00",
    87 => x"20",
    88 => x"51",
    89 => x"cf",
    90 => x"ff",
    91 => x"fa",
    92 => x"23",
    93 => x"fc",
    94 => x"00",
    95 => x"00",
    96 => x"00",
    97 => x"00",
    98 => x"00",
    99 => x"7f",
   100 => x"00",
   101 => x"52",
   102 => x"41",
   103 => x"fa",
   104 => x"00",
   105 => x"44",
   106 => x"61",
   107 => x"00",
   108 => x"06",
   109 => x"b8",
   110 => x"61",
   111 => x"00",
   112 => x"0a",
   113 => x"ea",
   114 => x"4a",
   115 => x"80",
   116 => x"67",
   117 => x"0a",
   118 => x"41",
   119 => x"fa",
   120 => x"00",
   121 => x"68",
   122 => x"61",
   123 => x"00",
   124 => x"06",
   125 => x"a8",
   126 => x"60",
   127 => x"fe",
   128 => x"41",
   129 => x"fa",
   130 => x"00",
   131 => x"47",
   132 => x"61",
   133 => x"00",
   134 => x"06",
   135 => x"9e",
   136 => x"61",
   137 => x"00",
   138 => x"02",
   139 => x"aa",
   140 => x"4b",
   141 => x"f9",
   142 => x"80",
   143 => x"00",
   144 => x"08",
   145 => x"00",
   146 => x"33",
   147 => x"fc",
   148 => x"00",
   149 => x"00",
   150 => x"00",
   151 => x"7f",
   152 => x"00",
   153 => x"0c",
   154 => x"30",
   155 => x"39",
   156 => x"81",
   157 => x"00",
   158 => x"00",
   159 => x"00",
   160 => x"08",
   161 => x"00",
   162 => x"00",
   163 => x"09",
   164 => x"67",
   165 => x"f4",
   166 => x"61",
   167 => x"00",
   168 => x"00",
   169 => x"80",
   170 => x"60",
   171 => x"ee",
   172 => x"43",
   173 => x"6f",
   174 => x"6e",
   175 => x"64",
   176 => x"75",
   177 => x"63",
   178 => x"74",
   179 => x"69",
   180 => x"6e",
   181 => x"67",
   182 => x"20",
   183 => x"73",
   184 => x"61",
   185 => x"6e",
   186 => x"69",
   187 => x"74",
   188 => x"79",
   189 => x"20",
   190 => x"63",
   191 => x"68",
   192 => x"65",
   193 => x"63",
   194 => x"6b",
   195 => x"2e",
   196 => x"2e",
   197 => x"2e",
   198 => x"0d",
   199 => x"0a",
   200 => x"00",
   201 => x"53",
   202 => x"61",
   203 => x"6e",
   204 => x"69",
   205 => x"74",
   206 => x"79",
   207 => x"20",
   208 => x"63",
   209 => x"68",
   210 => x"65",
   211 => x"63",
   212 => x"6b",
   213 => x"20",
   214 => x"70",
   215 => x"61",
   216 => x"73",
   217 => x"73",
   218 => x"65",
   219 => x"64",
   220 => x"2e",
   221 => x"0d",
   222 => x"0a",
   223 => x"00",
   224 => x"53",
   225 => x"61",
   226 => x"6e",
   227 => x"69",
   228 => x"74",
   229 => x"79",
   230 => x"20",
   231 => x"63",
   232 => x"68",
   233 => x"65",
   234 => x"63",
   235 => x"6b",
   236 => x"20",
   237 => x"66",
   238 => x"61",
   239 => x"69",
   240 => x"6c",
   241 => x"65",
   242 => x"64",
   243 => x"2e",
   244 => x"0d",
   245 => x"0a",
   246 => x"00",
   247 => x"00",
   248 => x"c0",
   249 => x"bc",
   250 => x"00",
   251 => x"00",
   252 => x"00",
   253 => x"df",
   254 => x"90",
   255 => x"3c",
   256 => x"00",
   257 => x"37",
   258 => x"6a",
   259 => x"04",
   260 => x"d0",
   261 => x"3c",
   262 => x"00",
   263 => x"27",
   264 => x"e9",
   265 => x"8e",
   266 => x"8c",
   267 => x"00",
   268 => x"20",
   269 => x"86",
   270 => x"4e",
   271 => x"75",
   272 => x"c0",
   273 => x"bc",
   274 => x"00",
   275 => x"00",
   276 => x"00",
   277 => x"df",
   278 => x"90",
   279 => x"3c",
   280 => x"00",
   281 => x"37",
   282 => x"6a",
   283 => x"04",
   284 => x"d0",
   285 => x"3c",
   286 => x"00",
   287 => x"27",
   288 => x"e9",
   289 => x"0f",
   290 => x"8e",
   291 => x"00",
   292 => x"10",
   293 => x"87",
   294 => x"4e",
   295 => x"75",
   296 => x"52",
   297 => x"79",
   298 => x"00",
   299 => x"7f",
   300 => x"00",
   301 => x"0c",
   302 => x"b0",
   303 => x"3c",
   304 => x"00",
   305 => x"53",
   306 => x"66",
   307 => x"2a",
   308 => x"33",
   309 => x"fc",
   310 => x"ff",
   311 => x"ff",
   312 => x"81",
   313 => x"00",
   314 => x"00",
   315 => x"06",
   316 => x"72",
   317 => x"00",
   318 => x"2e",
   319 => x"01",
   320 => x"2c",
   321 => x"01",
   322 => x"33",
   323 => x"c1",
   324 => x"00",
   325 => x"7f",
   326 => x"00",
   327 => x"0c",
   328 => x"23",
   329 => x"c1",
   330 => x"00",
   331 => x"7f",
   332 => x"00",
   333 => x"08",
   334 => x"23",
   335 => x"c1",
   336 => x"00",
   337 => x"7f",
   338 => x"00",
   339 => x"04",
   340 => x"23",
   341 => x"c1",
   342 => x"00",
   343 => x"7f",
   344 => x"00",
   345 => x"10",
   346 => x"60",
   347 => x"00",
   348 => x"01",
   349 => x"72",
   350 => x"2c",
   351 => x"39",
   352 => x"00",
   353 => x"7f",
   354 => x"00",
   355 => x"20",
   356 => x"2e",
   357 => x"39",
   358 => x"00",
   359 => x"7f",
   360 => x"00",
   361 => x"1c",
   362 => x"0c",
   363 => x"79",
   364 => x"00",
   365 => x"01",
   366 => x"00",
   367 => x"7f",
   368 => x"00",
   369 => x"0c",
   370 => x"66",
   371 => x"34",
   372 => x"33",
   373 => x"fc",
   374 => x"f0",
   375 => x"00",
   376 => x"81",
   377 => x"00",
   378 => x"00",
   379 => x"06",
   380 => x"41",
   381 => x"f9",
   382 => x"00",
   383 => x"7f",
   384 => x"00",
   385 => x"13",
   386 => x"61",
   387 => x"8c",
   388 => x"22",
   389 => x"39",
   390 => x"00",
   391 => x"7f",
   392 => x"00",
   393 => x"10",
   394 => x"b2",
   395 => x"bc",
   396 => x"00",
   397 => x"00",
   398 => x"00",
   399 => x"03",
   400 => x"6f",
   401 => x"08",
   402 => x"72",
   403 => x"0a",
   404 => x"92",
   405 => x"b9",
   406 => x"00",
   407 => x"7f",
   408 => x"00",
   409 => x"10",
   410 => x"52",
   411 => x"81",
   412 => x"e3",
   413 => x"89",
   414 => x"23",
   415 => x"c1",
   416 => x"00",
   417 => x"7f",
   418 => x"00",
   419 => x"14",
   420 => x"60",
   421 => x"00",
   422 => x"01",
   423 => x"28",
   424 => x"33",
   425 => x"f9",
   426 => x"00",
   427 => x"7f",
   428 => x"00",
   429 => x"12",
   430 => x"81",
   431 => x"00",
   432 => x"00",
   433 => x"06",
   434 => x"4a",
   435 => x"b9",
   436 => x"00",
   437 => x"7f",
   438 => x"00",
   439 => x"10",
   440 => x"67",
   441 => x"00",
   442 => x"01",
   443 => x"14",
   444 => x"0c",
   445 => x"b9",
   446 => x"00",
   447 => x"00",
   448 => x"00",
   449 => x"09",
   450 => x"00",
   451 => x"7f",
   452 => x"00",
   453 => x"10",
   454 => x"6e",
   455 => x"00",
   456 => x"00",
   457 => x"c0",
   458 => x"0c",
   459 => x"79",
   460 => x"00",
   461 => x"03",
   462 => x"00",
   463 => x"7f",
   464 => x"00",
   465 => x"0c",
   466 => x"6e",
   467 => x"16",
   468 => x"33",
   469 => x"fc",
   470 => x"0f",
   471 => x"00",
   472 => x"81",
   473 => x"00",
   474 => x"00",
   475 => x"06",
   476 => x"41",
   477 => x"f9",
   478 => x"00",
   479 => x"7f",
   480 => x"00",
   481 => x"07",
   482 => x"61",
   483 => x"00",
   484 => x"ff",
   485 => x"2c",
   486 => x"60",
   487 => x"00",
   488 => x"00",
   489 => x"e6",
   490 => x"22",
   491 => x"39",
   492 => x"00",
   493 => x"7f",
   494 => x"00",
   495 => x"14",
   496 => x"56",
   497 => x"41",
   498 => x"34",
   499 => x"39",
   500 => x"00",
   501 => x"7f",
   502 => x"00",
   503 => x"0c",
   504 => x"b4",
   505 => x"41",
   506 => x"6e",
   507 => x"20",
   508 => x"41",
   509 => x"f9",
   510 => x"00",
   511 => x"7f",
   512 => x"00",
   513 => x"08",
   514 => x"61",
   515 => x"00",
   516 => x"fe",
   517 => x"f4",
   518 => x"33",
   519 => x"f9",
   520 => x"00",
   521 => x"7f",
   522 => x"00",
   523 => x"0a",
   524 => x"81",
   525 => x"00",
   526 => x"00",
   527 => x"06",
   528 => x"33",
   529 => x"fc",
   530 => x"00",
   531 => x"01",
   532 => x"00",
   533 => x"7f",
   534 => x"00",
   535 => x"18",
   536 => x"60",
   537 => x"00",
   538 => x"00",
   539 => x"b4",
   540 => x"0c",
   541 => x"b9",
   542 => x"00",
   543 => x"00",
   544 => x"00",
   545 => x"03",
   546 => x"00",
   547 => x"7f",
   548 => x"00",
   549 => x"10",
   550 => x"6e",
   551 => x"60",
   552 => x"33",
   553 => x"fc",
   554 => x"00",
   555 => x"0f",
   556 => x"81",
   557 => x"00",
   558 => x"00",
   559 => x"06",
   560 => x"22",
   561 => x"39",
   562 => x"00",
   563 => x"7f",
   564 => x"00",
   565 => x"04",
   566 => x"e3",
   567 => x"89",
   568 => x"52",
   569 => x"81",
   570 => x"34",
   571 => x"39",
   572 => x"00",
   573 => x"7f",
   574 => x"00",
   575 => x"0c",
   576 => x"b4",
   577 => x"41",
   578 => x"6e",
   579 => x"2a",
   580 => x"20",
   581 => x"79",
   582 => x"00",
   583 => x"7f",
   584 => x"00",
   585 => x"08",
   586 => x"61",
   587 => x"00",
   588 => x"fe",
   589 => x"c4",
   590 => x"32",
   591 => x"39",
   592 => x"00",
   593 => x"7f",
   594 => x"00",
   595 => x"18",
   596 => x"53",
   597 => x"79",
   598 => x"00",
   599 => x"7f",
   600 => x"00",
   601 => x"18",
   602 => x"53",
   603 => x"41",
   604 => x"6a",
   605 => x"70",
   606 => x"52",
   607 => x"b9",
   608 => x"00",
   609 => x"7f",
   610 => x"00",
   611 => x"08",
   612 => x"33",
   613 => x"fc",
   614 => x"00",
   615 => x"01",
   616 => x"00",
   617 => x"7f",
   618 => x"00",
   619 => x"18",
   620 => x"60",
   621 => x"60",
   622 => x"30",
   623 => x"39",
   624 => x"00",
   625 => x"7f",
   626 => x"00",
   627 => x"18",
   628 => x"52",
   629 => x"40",
   630 => x"c0",
   631 => x"7c",
   632 => x"00",
   633 => x"01",
   634 => x"67",
   635 => x"52",
   636 => x"20",
   637 => x"79",
   638 => x"00",
   639 => x"7f",
   640 => x"00",
   641 => x"08",
   642 => x"e5",
   643 => x"88",
   644 => x"e1",
   645 => x"2f",
   646 => x"10",
   647 => x"87",
   648 => x"33",
   649 => x"fc",
   650 => x"f0",
   651 => x"f0",
   652 => x"81",
   653 => x"00",
   654 => x"00",
   655 => x"06",
   656 => x"0c",
   657 => x"b9",
   658 => x"00",
   659 => x"00",
   660 => x"00",
   661 => x"07",
   662 => x"00",
   663 => x"7f",
   664 => x"00",
   665 => x"10",
   666 => x"6d",
   667 => x"32",
   668 => x"33",
   669 => x"fc",
   670 => x"f0",
   671 => x"0f",
   672 => x"81",
   673 => x"00",
   674 => x"00",
   675 => x"06",
   676 => x"0c",
   677 => x"b9",
   678 => x"00",
   679 => x"00",
   680 => x"00",
   681 => x"09",
   682 => x"00",
   683 => x"7f",
   684 => x"00",
   685 => x"10",
   686 => x"6e",
   687 => x"1e",
   688 => x"33",
   689 => x"fc",
   690 => x"ff",
   691 => x"f0",
   692 => x"81",
   693 => x"00",
   694 => x"00",
   695 => x"06",
   696 => x"41",
   697 => x"fa",
   698 => x"00",
   699 => x"22",
   700 => x"61",
   701 => x"56",
   702 => x"2e",
   703 => x"b9",
   704 => x"00",
   705 => x"7f",
   706 => x"00",
   707 => x"08",
   708 => x"08",
   709 => x"b9",
   710 => x"00",
   711 => x"00",
   712 => x"81",
   713 => x"00",
   714 => x"00",
   715 => x"04",
   716 => x"4e",
   717 => x"75",
   718 => x"23",
   719 => x"c6",
   720 => x"00",
   721 => x"7f",
   722 => x"00",
   723 => x"20",
   724 => x"23",
   725 => x"c7",
   726 => x"00",
   727 => x"7f",
   728 => x"00",
   729 => x"1c",
   730 => x"4e",
   731 => x"75",
   732 => x"46",
   733 => x"69",
   734 => x"72",
   735 => x"6d",
   736 => x"77",
   737 => x"61",
   738 => x"72",
   739 => x"65",
   740 => x"20",
   741 => x"72",
   742 => x"65",
   743 => x"63",
   744 => x"65",
   745 => x"69",
   746 => x"76",
   747 => x"65",
   748 => x"64",
   749 => x"20",
   750 => x"2d",
   751 => x"20",
   752 => x"6c",
   753 => x"61",
   754 => x"75",
   755 => x"6e",
   756 => x"63",
   757 => x"68",
   758 => x"69",
   759 => x"6e",
   760 => x"67",
   761 => x"0d",
   762 => x"0a",
   763 => x"00",
   764 => x"48",
   765 => x"40",
   766 => x"30",
   767 => x"39",
   768 => x"81",
   769 => x"00",
   770 => x"00",
   771 => x"00",
   772 => x"08",
   773 => x"00",
   774 => x"00",
   775 => x"08",
   776 => x"67",
   777 => x"f4",
   778 => x"48",
   779 => x"40",
   780 => x"33",
   781 => x"c0",
   782 => x"81",
   783 => x"00",
   784 => x"00",
   785 => x"00",
   786 => x"4e",
   787 => x"75",
   788 => x"2f",
   789 => x"00",
   790 => x"70",
   791 => x"00",
   792 => x"30",
   793 => x"39",
   794 => x"81",
   795 => x"00",
   796 => x"00",
   797 => x"00",
   798 => x"08",
   799 => x"00",
   800 => x"00",
   801 => x"08",
   802 => x"67",
   803 => x"f4",
   804 => x"10",
   805 => x"18",
   806 => x"67",
   807 => x"08",
   808 => x"33",
   809 => x"c0",
   810 => x"81",
   811 => x"00",
   812 => x"00",
   813 => x"00",
   814 => x"60",
   815 => x"e8",
   816 => x"20",
   817 => x"1f",
   818 => x"4e",
   819 => x"75",
   820 => x"33",
   821 => x"fc",
   822 => x"00",
   823 => x"01",
   824 => x"81",
   825 => x"00",
   826 => x"00",
   827 => x"06",
   828 => x"41",
   829 => x"fa",
   830 => x"01",
   831 => x"fa",
   832 => x"61",
   833 => x"00",
   834 => x"03",
   835 => x"e2",
   836 => x"61",
   837 => x"00",
   838 => x"02",
   839 => x"60",
   840 => x"66",
   841 => x"5c",
   842 => x"33",
   843 => x"fc",
   844 => x"00",
   845 => x"02",
   846 => x"81",
   847 => x"00",
   848 => x"00",
   849 => x"06",
   850 => x"33",
   851 => x"fc",
   852 => x"00",
   853 => x"40",
   854 => x"00",
   855 => x"7f",
   856 => x"00",
   857 => x"26",
   858 => x"61",
   859 => x"00",
   860 => x"04",
   861 => x"8a",
   862 => x"67",
   863 => x"0c",
   864 => x"42",
   865 => x"79",
   866 => x"00",
   867 => x"7f",
   868 => x"00",
   869 => x"26",
   870 => x"61",
   871 => x"00",
   872 => x"04",
   873 => x"7e",
   874 => x"66",
   875 => x"28",
   876 => x"33",
   877 => x"fc",
   878 => x"00",
   879 => x"03",
   880 => x"81",
   881 => x"00",
   882 => x"00",
   883 => x"06",
   884 => x"61",
   885 => x"00",
   886 => x"05",
   887 => x"f8",
   888 => x"43",
   889 => x"fa",
   890 => x"00",
   891 => x"57",
   892 => x"61",
   893 => x"00",
   894 => x"06",
   895 => x"48",
   896 => x"67",
   897 => x"12",
   898 => x"41",
   899 => x"fa",
   900 => x"00",
   901 => x"47",
   902 => x"61",
   903 => x"00",
   904 => x"03",
   905 => x"9c",
   906 => x"30",
   907 => x"7c",
   908 => x"20",
   909 => x"00",
   910 => x"61",
   911 => x"00",
   912 => x"04",
   913 => x"02",
   914 => x"4e",
   915 => x"75",
   916 => x"33",
   917 => x"fc",
   918 => x"f0",
   919 => x"03",
   920 => x"81",
   921 => x"00",
   922 => x"00",
   923 => x"06",
   924 => x"41",
   925 => x"fa",
   926 => x"00",
   927 => x"29",
   928 => x"61",
   929 => x"00",
   930 => x"03",
   931 => x"82",
   932 => x"4e",
   933 => x"75",
   934 => x"33",
   935 => x"fc",
   936 => x"f0",
   937 => x"02",
   938 => x"81",
   939 => x"00",
   940 => x"00",
   941 => x"06",
   942 => x"41",
   943 => x"fa",
   944 => x"00",
   945 => x"08",
   946 => x"61",
   947 => x"00",
   948 => x"03",
   949 => x"70",
   950 => x"4e",
   951 => x"75",
   952 => x"53",
   953 => x"44",
   954 => x"20",
   955 => x"69",
   956 => x"6e",
   957 => x"69",
   958 => x"74",
   959 => x"20",
   960 => x"66",
   961 => x"61",
   962 => x"69",
   963 => x"6c",
   964 => x"65",
   965 => x"64",
   966 => x"00",
   967 => x"6e",
   968 => x"6f",
   969 => x"74",
   970 => x"20",
   971 => x"66",
   972 => x"6f",
   973 => x"75",
   974 => x"6e",
   975 => x"64",
   976 => x"20",
   977 => x"42",
   978 => x"4f",
   979 => x"4f",
   980 => x"54",
   981 => x"20",
   982 => x"20",
   983 => x"20",
   984 => x"20",
   985 => x"53",
   986 => x"52",
   987 => x"45",
   988 => x"00",
   989 => x"00",
   990 => x"33",
   991 => x"fc",
   992 => x"01",
   993 => x"00",
   994 => x"81",
   995 => x"00",
   996 => x"00",
   997 => x"06",
   998 => x"41",
   999 => x"f9",
  1000 => x"00",
  1001 => x"7f",
  1002 => x"00",
  1003 => x"56",
  1004 => x"61",
  1005 => x"00",
  1006 => x"00",
  1007 => x"c4",
  1008 => x"66",
  1009 => x"68",
  1010 => x"33",
  1011 => x"fc",
  1012 => x"01",
  1013 => x"01",
  1014 => x"81",
  1015 => x"00",
  1016 => x"00",
  1017 => x"06",
  1018 => x"32",
  1019 => x"3c",
  1020 => x"4e",
  1021 => x"20",
  1022 => x"53",
  1023 => x"41",
  1024 => x"67",
  1025 => x"44",
  1026 => x"33",
  1027 => x"fc",
  1028 => x"01",
  1029 => x"02",
  1030 => x"81",
  1031 => x"00",
  1032 => x"00",
  1033 => x"06",
  1034 => x"33",
  1035 => x"7c",
  1036 => x"00",
  1037 => x"ff",
  1038 => x"00",
  1039 => x"24",
  1040 => x"30",
  1041 => x"29",
  1042 => x"00",
  1043 => x"24",
  1044 => x"b0",
  1045 => x"3c",
  1046 => x"00",
  1047 => x"fe",
  1048 => x"66",
  1049 => x"e4",
  1050 => x"30",
  1051 => x"29",
  1052 => x"01",
  1053 => x"00",
  1054 => x"32",
  1055 => x"3c",
  1056 => x"00",
  1057 => x"7f",
  1058 => x"20",
  1059 => x"29",
  1060 => x"01",
  1061 => x"00",
  1062 => x"20",
  1063 => x"c0",
  1064 => x"51",
  1065 => x"c9",
  1066 => x"ff",
  1067 => x"f8",
  1068 => x"30",
  1069 => x"29",
  1070 => x"00",
  1071 => x"24",
  1072 => x"33",
  1073 => x"7c",
  1074 => x"00",
  1075 => x"00",
  1076 => x"00",
  1077 => x"22",
  1078 => x"33",
  1079 => x"fc",
  1080 => x"01",
  1081 => x"03",
  1082 => x"81",
  1083 => x"00",
  1084 => x"00",
  1085 => x"06",
  1086 => x"41",
  1087 => x"e8",
  1088 => x"fe",
  1089 => x"00",
  1090 => x"70",
  1091 => x"00",
  1092 => x"4e",
  1093 => x"75",
  1094 => x"33",
  1095 => x"fc",
  1096 => x"f1",
  1097 => x"02",
  1098 => x"81",
  1099 => x"00",
  1100 => x"00",
  1101 => x"06",
  1102 => x"41",
  1103 => x"fa",
  1104 => x"01",
  1105 => x"38",
  1106 => x"61",
  1107 => x"00",
  1108 => x"02",
  1109 => x"d0",
  1110 => x"70",
  1111 => x"fe",
  1112 => x"4e",
  1113 => x"75",
  1114 => x"33",
  1115 => x"fc",
  1116 => x"f1",
  1117 => x"03",
  1118 => x"81",
  1119 => x"00",
  1120 => x"00",
  1121 => x"06",
  1122 => x"41",
  1123 => x"fa",
  1124 => x"01",
  1125 => x"0c",
  1126 => x"61",
  1127 => x"00",
  1128 => x"02",
  1129 => x"bc",
  1130 => x"70",
  1131 => x"ff",
  1132 => x"4e",
  1133 => x"75",
  1134 => x"22",
  1135 => x"3c",
  1136 => x"00",
  1137 => x"95",
  1138 => x"00",
  1139 => x"40",
  1140 => x"70",
  1141 => x"00",
  1142 => x"60",
  1143 => x"40",
  1144 => x"22",
  1145 => x"3c",
  1146 => x"00",
  1147 => x"ff",
  1148 => x"00",
  1149 => x"41",
  1150 => x"70",
  1151 => x"00",
  1152 => x"60",
  1153 => x"36",
  1154 => x"22",
  1155 => x"3c",
  1156 => x"00",
  1157 => x"87",
  1158 => x"00",
  1159 => x"48",
  1160 => x"20",
  1161 => x"3c",
  1162 => x"00",
  1163 => x"00",
  1164 => x"01",
  1165 => x"aa",
  1166 => x"60",
  1167 => x"28",
  1168 => x"22",
  1169 => x"3c",
  1170 => x"00",
  1171 => x"87",
  1172 => x"00",
  1173 => x"69",
  1174 => x"20",
  1175 => x"3c",
  1176 => x"40",
  1177 => x"00",
  1178 => x"00",
  1179 => x"00",
  1180 => x"60",
  1181 => x"1a",
  1182 => x"22",
  1183 => x"3c",
  1184 => x"00",
  1185 => x"ff",
  1186 => x"00",
  1187 => x"77",
  1188 => x"70",
  1189 => x"00",
  1190 => x"60",
  1191 => x"10",
  1192 => x"22",
  1193 => x"3c",
  1194 => x"00",
  1195 => x"ff",
  1196 => x"00",
  1197 => x"7a",
  1198 => x"70",
  1199 => x"00",
  1200 => x"60",
  1201 => x"06",
  1202 => x"22",
  1203 => x"3c",
  1204 => x"00",
  1205 => x"ff",
  1206 => x"00",
  1207 => x"51",
  1208 => x"43",
  1209 => x"f9",
  1210 => x"81",
  1211 => x"00",
  1212 => x"00",
  1213 => x"00",
  1214 => x"33",
  1215 => x"7c",
  1216 => x"00",
  1217 => x"ff",
  1218 => x"00",
  1219 => x"24",
  1220 => x"3f",
  1221 => x"69",
  1222 => x"00",
  1223 => x"24",
  1224 => x"ff",
  1225 => x"fe",
  1226 => x"33",
  1227 => x"7c",
  1228 => x"00",
  1229 => x"01",
  1230 => x"00",
  1231 => x"22",
  1232 => x"33",
  1233 => x"7c",
  1234 => x"00",
  1235 => x"ff",
  1236 => x"00",
  1237 => x"24",
  1238 => x"33",
  1239 => x"41",
  1240 => x"00",
  1241 => x"24",
  1242 => x"48",
  1243 => x"41",
  1244 => x"4a",
  1245 => x"79",
  1246 => x"00",
  1247 => x"7f",
  1248 => x"00",
  1249 => x"24",
  1250 => x"67",
  1251 => x"16",
  1252 => x"e1",
  1253 => x"98",
  1254 => x"33",
  1255 => x"40",
  1256 => x"00",
  1257 => x"24",
  1258 => x"e1",
  1259 => x"98",
  1260 => x"33",
  1261 => x"40",
  1262 => x"00",
  1263 => x"24",
  1264 => x"e1",
  1265 => x"98",
  1266 => x"33",
  1267 => x"40",
  1268 => x"00",
  1269 => x"24",
  1270 => x"e1",
  1271 => x"98",
  1272 => x"60",
  1273 => x"18",
  1274 => x"d0",
  1275 => x"80",
  1276 => x"48",
  1277 => x"40",
  1278 => x"33",
  1279 => x"40",
  1280 => x"00",
  1281 => x"24",
  1282 => x"48",
  1283 => x"40",
  1284 => x"e1",
  1285 => x"58",
  1286 => x"33",
  1287 => x"40",
  1288 => x"00",
  1289 => x"24",
  1290 => x"e1",
  1291 => x"58",
  1292 => x"33",
  1293 => x"40",
  1294 => x"00",
  1295 => x"24",
  1296 => x"70",
  1297 => x"00",
  1298 => x"33",
  1299 => x"40",
  1300 => x"00",
  1301 => x"24",
  1302 => x"33",
  1303 => x"41",
  1304 => x"00",
  1305 => x"24",
  1306 => x"22",
  1307 => x"3c",
  1308 => x"00",
  1309 => x"00",
  1310 => x"01",
  1311 => x"90",
  1312 => x"53",
  1313 => x"81",
  1314 => x"67",
  1315 => x"10",
  1316 => x"33",
  1317 => x"7c",
  1318 => x"00",
  1319 => x"ff",
  1320 => x"00",
  1321 => x"24",
  1322 => x"30",
  1323 => x"29",
  1324 => x"00",
  1325 => x"24",
  1326 => x"b0",
  1327 => x"3c",
  1328 => x"00",
  1329 => x"ff",
  1330 => x"67",
  1331 => x"ec",
  1332 => x"80",
  1333 => x"00",
  1334 => x"4e",
  1335 => x"75",
  1336 => x"53",
  1337 => x"74",
  1338 => x"61",
  1339 => x"72",
  1340 => x"74",
  1341 => x"20",
  1342 => x"49",
  1343 => x"6e",
  1344 => x"69",
  1345 => x"74",
  1346 => x"0d",
  1347 => x"0a",
  1348 => x"00",
  1349 => x"49",
  1350 => x"6e",
  1351 => x"69",
  1352 => x"74",
  1353 => x"20",
  1354 => x"64",
  1355 => x"6f",
  1356 => x"6e",
  1357 => x"65",
  1358 => x"0d",
  1359 => x"0a",
  1360 => x"00",
  1361 => x"49",
  1362 => x"6e",
  1363 => x"69",
  1364 => x"74",
  1365 => x"20",
  1366 => x"66",
  1367 => x"61",
  1368 => x"69",
  1369 => x"6c",
  1370 => x"75",
  1371 => x"72",
  1372 => x"65",
  1373 => x"0d",
  1374 => x"0a",
  1375 => x"00",
  1376 => x"52",
  1377 => x"65",
  1378 => x"73",
  1379 => x"65",
  1380 => x"74",
  1381 => x"20",
  1382 => x"66",
  1383 => x"61",
  1384 => x"69",
  1385 => x"6c",
  1386 => x"75",
  1387 => x"72",
  1388 => x"65",
  1389 => x"0d",
  1390 => x"0a",
  1391 => x"00",
  1392 => x"43",
  1393 => x"6f",
  1394 => x"6d",
  1395 => x"6d",
  1396 => x"61",
  1397 => x"6e",
  1398 => x"64",
  1399 => x"20",
  1400 => x"54",
  1401 => x"69",
  1402 => x"6d",
  1403 => x"65",
  1404 => x"6f",
  1405 => x"75",
  1406 => x"74",
  1407 => x"5f",
  1408 => x"45",
  1409 => x"72",
  1410 => x"72",
  1411 => x"6f",
  1412 => x"72",
  1413 => x"0d",
  1414 => x"0a",
  1415 => x"00",
  1416 => x"54",
  1417 => x"69",
  1418 => x"6d",
  1419 => x"65",
  1420 => x"6f",
  1421 => x"75",
  1422 => x"74",
  1423 => x"5f",
  1424 => x"45",
  1425 => x"72",
  1426 => x"72",
  1427 => x"6f",
  1428 => x"72",
  1429 => x"0d",
  1430 => x"0a",
  1431 => x"00",
  1432 => x"53",
  1433 => x"44",
  1434 => x"48",
  1435 => x"43",
  1436 => x"20",
  1437 => x"66",
  1438 => x"6f",
  1439 => x"75",
  1440 => x"6e",
  1441 => x"64",
  1442 => x"20",
  1443 => x"0d",
  1444 => x"0a",
  1445 => x"00",
  1446 => x"33",
  1447 => x"fc",
  1448 => x"ff",
  1449 => x"ff",
  1450 => x"00",
  1451 => x"7f",
  1452 => x"00",
  1453 => x"24",
  1454 => x"43",
  1455 => x"f9",
  1456 => x"81",
  1457 => x"00",
  1458 => x"00",
  1459 => x"00",
  1460 => x"33",
  1461 => x"7c",
  1462 => x"00",
  1463 => x"00",
  1464 => x"00",
  1465 => x"22",
  1466 => x"33",
  1467 => x"7c",
  1468 => x"00",
  1469 => x"96",
  1470 => x"00",
  1471 => x"1e",
  1472 => x"32",
  1473 => x"3c",
  1474 => x"00",
  1475 => x"c8",
  1476 => x"43",
  1477 => x"e9",
  1478 => x"00",
  1479 => x"20",
  1480 => x"33",
  1481 => x"7c",
  1482 => x"00",
  1483 => x"ff",
  1484 => x"00",
  1485 => x"24",
  1486 => x"51",
  1487 => x"c9",
  1488 => x"ff",
  1489 => x"f8",
  1490 => x"34",
  1491 => x"3c",
  1492 => x"00",
  1493 => x"32",
  1494 => x"61",
  1495 => x"00",
  1496 => x"fe",
  1497 => x"96",
  1498 => x"3f",
  1499 => x"69",
  1500 => x"00",
  1501 => x"24",
  1502 => x"ff",
  1503 => x"fe",
  1504 => x"33",
  1505 => x"7c",
  1506 => x"00",
  1507 => x"00",
  1508 => x"00",
  1509 => x"22",
  1510 => x"b0",
  1511 => x"3c",
  1512 => x"00",
  1513 => x"01",
  1514 => x"67",
  1515 => x"12",
  1516 => x"51",
  1517 => x"ca",
  1518 => x"ff",
  1519 => x"e8",
  1520 => x"48",
  1521 => x"7a",
  1522 => x"ff",
  1523 => x"6e",
  1524 => x"61",
  1525 => x"00",
  1526 => x"01",
  1527 => x"22",
  1528 => x"58",
  1529 => x"8f",
  1530 => x"70",
  1531 => x"ff",
  1532 => x"4e",
  1533 => x"75",
  1534 => x"22",
  1535 => x"3c",
  1536 => x"00",
  1537 => x"00",
  1538 => x"20",
  1539 => x"00",
  1540 => x"33",
  1541 => x"7c",
  1542 => x"00",
  1543 => x"ff",
  1544 => x"00",
  1545 => x"24",
  1546 => x"53",
  1547 => x"81",
  1548 => x"66",
  1549 => x"f6",
  1550 => x"61",
  1551 => x"00",
  1552 => x"fe",
  1553 => x"72",
  1554 => x"b0",
  1555 => x"3c",
  1556 => x"00",
  1557 => x"01",
  1558 => x"66",
  1559 => x"00",
  1560 => x"00",
  1561 => x"9e",
  1562 => x"33",
  1563 => x"7c",
  1564 => x"00",
  1565 => x"ff",
  1566 => x"00",
  1567 => x"24",
  1568 => x"33",
  1569 => x"7c",
  1570 => x"00",
  1571 => x"ff",
  1572 => x"00",
  1573 => x"24",
  1574 => x"33",
  1575 => x"7c",
  1576 => x"00",
  1577 => x"ff",
  1578 => x"00",
  1579 => x"24",
  1580 => x"30",
  1581 => x"29",
  1582 => x"00",
  1583 => x"24",
  1584 => x"0c",
  1585 => x"00",
  1586 => x"00",
  1587 => x"01",
  1588 => x"66",
  1589 => x"00",
  1590 => x"00",
  1591 => x"80",
  1592 => x"33",
  1593 => x"7c",
  1594 => x"00",
  1595 => x"ff",
  1596 => x"00",
  1597 => x"24",
  1598 => x"30",
  1599 => x"29",
  1600 => x"00",
  1601 => x"24",
  1602 => x"0c",
  1603 => x"00",
  1604 => x"00",
  1605 => x"aa",
  1606 => x"66",
  1607 => x"6e",
  1608 => x"3f",
  1609 => x"69",
  1610 => x"00",
  1611 => x"24",
  1612 => x"ff",
  1613 => x"fe",
  1614 => x"33",
  1615 => x"7c",
  1616 => x"00",
  1617 => x"00",
  1618 => x"00",
  1619 => x"22",
  1620 => x"48",
  1621 => x"7a",
  1622 => x"ff",
  1623 => x"42",
  1624 => x"61",
  1625 => x"00",
  1626 => x"00",
  1627 => x"be",
  1628 => x"58",
  1629 => x"8f",
  1630 => x"34",
  1631 => x"3c",
  1632 => x"00",
  1633 => x"32",
  1634 => x"53",
  1635 => x"42",
  1636 => x"67",
  1637 => x"50",
  1638 => x"32",
  1639 => x"3c",
  1640 => x"07",
  1641 => x"d0",
  1642 => x"33",
  1643 => x"7c",
  1644 => x"00",
  1645 => x"ff",
  1646 => x"00",
  1647 => x"24",
  1648 => x"51",
  1649 => x"c9",
  1650 => x"ff",
  1651 => x"f8",
  1652 => x"61",
  1653 => x"00",
  1654 => x"fe",
  1655 => x"28",
  1656 => x"b0",
  1657 => x"3c",
  1658 => x"00",
  1659 => x"01",
  1660 => x"66",
  1661 => x"e4",
  1662 => x"61",
  1663 => x"00",
  1664 => x"fe",
  1665 => x"10",
  1666 => x"66",
  1667 => x"de",
  1668 => x"61",
  1669 => x"00",
  1670 => x"fe",
  1671 => x"22",
  1672 => x"66",
  1673 => x"d8",
  1674 => x"33",
  1675 => x"7c",
  1676 => x"00",
  1677 => x"ff",
  1678 => x"00",
  1679 => x"24",
  1680 => x"30",
  1681 => x"29",
  1682 => x"00",
  1683 => x"24",
  1684 => x"c0",
  1685 => x"3c",
  1686 => x"00",
  1687 => x"40",
  1688 => x"66",
  1689 => x"08",
  1690 => x"33",
  1691 => x"fc",
  1692 => x"00",
  1693 => x"00",
  1694 => x"00",
  1695 => x"7f",
  1696 => x"00",
  1697 => x"24",
  1698 => x"33",
  1699 => x"7c",
  1700 => x"00",
  1701 => x"ff",
  1702 => x"00",
  1703 => x"24",
  1704 => x"33",
  1705 => x"7c",
  1706 => x"00",
  1707 => x"ff",
  1708 => x"00",
  1709 => x"24",
  1710 => x"33",
  1711 => x"7c",
  1712 => x"00",
  1713 => x"ff",
  1714 => x"00",
  1715 => x"24",
  1716 => x"60",
  1717 => x"3c",
  1718 => x"33",
  1719 => x"fc",
  1720 => x"00",
  1721 => x"00",
  1722 => x"00",
  1723 => x"7f",
  1724 => x"00",
  1725 => x"24",
  1726 => x"34",
  1727 => x"3c",
  1728 => x"00",
  1729 => x"0a",
  1730 => x"32",
  1731 => x"3c",
  1732 => x"07",
  1733 => x"d0",
  1734 => x"33",
  1735 => x"7c",
  1736 => x"00",
  1737 => x"ff",
  1738 => x"00",
  1739 => x"24",
  1740 => x"51",
  1741 => x"c9",
  1742 => x"ff",
  1743 => x"f8",
  1744 => x"61",
  1745 => x"00",
  1746 => x"fd",
  1747 => x"a6",
  1748 => x"67",
  1749 => x"1c",
  1750 => x"3f",
  1751 => x"69",
  1752 => x"00",
  1753 => x"24",
  1754 => x"ff",
  1755 => x"fe",
  1756 => x"33",
  1757 => x"7c",
  1758 => x"00",
  1759 => x"00",
  1760 => x"00",
  1761 => x"22",
  1762 => x"51",
  1763 => x"ca",
  1764 => x"ff",
  1765 => x"de",
  1766 => x"48",
  1767 => x"7a",
  1768 => x"fe",
  1769 => x"69",
  1770 => x"61",
  1771 => x"2c",
  1772 => x"58",
  1773 => x"8f",
  1774 => x"70",
  1775 => x"ff",
  1776 => x"4e",
  1777 => x"75",
  1778 => x"3f",
  1779 => x"69",
  1780 => x"00",
  1781 => x"24",
  1782 => x"ff",
  1783 => x"fe",
  1784 => x"33",
  1785 => x"7c",
  1786 => x"00",
  1787 => x"00",
  1788 => x"00",
  1789 => x"22",
  1790 => x"33",
  1791 => x"69",
  1792 => x"00",
  1793 => x"2c",
  1794 => x"00",
  1795 => x"1e",
  1796 => x"48",
  1797 => x"7a",
  1798 => x"fe",
  1799 => x"3f",
  1800 => x"61",
  1801 => x"0e",
  1802 => x"58",
  1803 => x"8f",
  1804 => x"33",
  1805 => x"fc",
  1806 => x"ff",
  1807 => x"ff",
  1808 => x"81",
  1809 => x"00",
  1810 => x"00",
  1811 => x"06",
  1812 => x"70",
  1813 => x"00",
  1814 => x"4e",
  1815 => x"75",
  1816 => x"2f",
  1817 => x"08",
  1818 => x"20",
  1819 => x"6f",
  1820 => x"00",
  1821 => x"08",
  1822 => x"61",
  1823 => x"04",
  1824 => x"20",
  1825 => x"5f",
  1826 => x"4e",
  1827 => x"75",
  1828 => x"48",
  1829 => x"e7",
  1830 => x"00",
  1831 => x"c0",
  1832 => x"22",
  1833 => x"39",
  1834 => x"00",
  1835 => x"7f",
  1836 => x"00",
  1837 => x"52",
  1838 => x"43",
  1839 => x"f9",
  1840 => x"80",
  1841 => x"00",
  1842 => x"08",
  1843 => x"00",
  1844 => x"10",
  1845 => x"18",
  1846 => x"67",
  1847 => x"08",
  1848 => x"13",
  1849 => x"80",
  1850 => x"10",
  1851 => x"00",
  1852 => x"52",
  1853 => x"41",
  1854 => x"60",
  1855 => x"f4",
  1856 => x"06",
  1857 => x"b9",
  1858 => x"00",
  1859 => x"00",
  1860 => x"00",
  1861 => x"4c",
  1862 => x"00",
  1863 => x"7f",
  1864 => x"00",
  1865 => x"52",
  1866 => x"4c",
  1867 => x"df",
  1868 => x"03",
  1869 => x"00",
  1870 => x"4e",
  1871 => x"75",
  1872 => x"4a",
  1873 => x"79",
  1874 => x"00",
  1875 => x"7f",
  1876 => x"00",
  1877 => x"24",
  1878 => x"67",
  1879 => x"1e",
  1880 => x"41",
  1881 => x"fa",
  1882 => x"00",
  1883 => x"08",
  1884 => x"48",
  1885 => x"7a",
  1886 => x"00",
  1887 => x"34",
  1888 => x"60",
  1889 => x"c2",
  1890 => x"53",
  1891 => x"44",
  1892 => x"48",
  1893 => x"43",
  1894 => x"20",
  1895 => x"66",
  1896 => x"6c",
  1897 => x"61",
  1898 => x"67",
  1899 => x"20",
  1900 => x"73",
  1901 => x"74",
  1902 => x"69",
  1903 => x"6c",
  1904 => x"6c",
  1905 => x"20",
  1906 => x"73",
  1907 => x"65",
  1908 => x"74",
  1909 => x"00",
  1910 => x"41",
  1911 => x"fa",
  1912 => x"00",
  1913 => x"08",
  1914 => x"48",
  1915 => x"7a",
  1916 => x"00",
  1917 => x"16",
  1918 => x"60",
  1919 => x"a4",
  1920 => x"53",
  1921 => x"44",
  1922 => x"48",
  1923 => x"43",
  1924 => x"20",
  1925 => x"66",
  1926 => x"6c",
  1927 => x"61",
  1928 => x"67",
  1929 => x"20",
  1930 => x"63",
  1931 => x"6c",
  1932 => x"65",
  1933 => x"61",
  1934 => x"72",
  1935 => x"65",
  1936 => x"64",
  1937 => x"00",
  1938 => x"61",
  1939 => x"00",
  1940 => x"02",
  1941 => x"0a",
  1942 => x"61",
  1943 => x"00",
  1944 => x"fc",
  1945 => x"46",
  1946 => x"66",
  1947 => x"46",
  1948 => x"2e",
  1949 => x"3c",
  1950 => x"00",
  1951 => x"00",
  1952 => x"01",
  1953 => x"ff",
  1954 => x"41",
  1955 => x"f9",
  1956 => x"00",
  1957 => x"7f",
  1958 => x"00",
  1959 => x"56",
  1960 => x"43",
  1961 => x"f9",
  1962 => x"80",
  1963 => x"00",
  1964 => x"08",
  1965 => x"00",
  1966 => x"10",
  1967 => x"18",
  1968 => x"12",
  1969 => x"c0",
  1970 => x"48",
  1971 => x"e7",
  1972 => x"01",
  1973 => x"c0",
  1974 => x"61",
  1975 => x"00",
  1976 => x"f9",
  1977 => x"70",
  1978 => x"4c",
  1979 => x"df",
  1980 => x"03",
  1981 => x"80",
  1982 => x"51",
  1983 => x"cf",
  1984 => x"ff",
  1985 => x"ee",
  1986 => x"20",
  1987 => x"39",
  1988 => x"00",
  1989 => x"7f",
  1990 => x"00",
  1991 => x"38",
  1992 => x"52",
  1993 => x"80",
  1994 => x"23",
  1995 => x"c0",
  1996 => x"00",
  1997 => x"7f",
  1998 => x"00",
  1999 => x"38",
  2000 => x"53",
  2001 => x"79",
  2002 => x"00",
  2003 => x"7f",
  2004 => x"00",
  2005 => x"36",
  2006 => x"66",
  2007 => x"be",
  2008 => x"61",
  2009 => x"00",
  2010 => x"02",
  2011 => x"7a",
  2012 => x"66",
  2013 => x"b4",
  2014 => x"20",
  2015 => x"08",
  2016 => x"4e",
  2017 => x"75",
  2018 => x"70",
  2019 => x"00",
  2020 => x"4e",
  2021 => x"75",
  2022 => x"33",
  2023 => x"fc",
  2024 => x"02",
  2025 => x"01",
  2026 => x"81",
  2027 => x"00",
  2028 => x"00",
  2029 => x"06",
  2030 => x"70",
  2031 => x"00",
  2032 => x"23",
  2033 => x"c0",
  2034 => x"00",
  2035 => x"7f",
  2036 => x"00",
  2037 => x"3e",
  2038 => x"33",
  2039 => x"fc",
  2040 => x"02",
  2041 => x"11",
  2042 => x"81",
  2043 => x"00",
  2044 => x"00",
  2045 => x"06",
  2046 => x"61",
  2047 => x"00",
  2048 => x"fb",
  2049 => x"de",
  2050 => x"66",
  2051 => x"5c",
  2052 => x"33",
  2053 => x"fc",
  2054 => x"02",
  2055 => x"02",
  2056 => x"81",
  2057 => x"00",
  2058 => x"00",
  2059 => x"06",
  2060 => x"0c",
  2061 => x"28",
  2062 => x"00",
  2063 => x"55",
  2064 => x"01",
  2065 => x"fe",
  2066 => x"66",
  2067 => x"4c",
  2068 => x"0c",
  2069 => x"28",
  2070 => x"00",
  2071 => x"aa",
  2072 => x"01",
  2073 => x"ff",
  2074 => x"66",
  2075 => x"44",
  2076 => x"30",
  2077 => x"39",
  2078 => x"00",
  2079 => x"7f",
  2080 => x"00",
  2081 => x"26",
  2082 => x"c0",
  2083 => x"7c",
  2084 => x"00",
  2085 => x"70",
  2086 => x"b0",
  2087 => x"7c",
  2088 => x"00",
  2089 => x"40",
  2090 => x"64",
  2091 => x"40",
  2092 => x"43",
  2093 => x"e8",
  2094 => x"01",
  2095 => x"be",
  2096 => x"d2",
  2097 => x"c0",
  2098 => x"33",
  2099 => x"fc",
  2100 => x"02",
  2101 => x"03",
  2102 => x"81",
  2103 => x"00",
  2104 => x"00",
  2105 => x"06",
  2106 => x"20",
  2107 => x"29",
  2108 => x"00",
  2109 => x"08",
  2110 => x"e0",
  2111 => x"58",
  2112 => x"48",
  2113 => x"40",
  2114 => x"e0",
  2115 => x"58",
  2116 => x"23",
  2117 => x"c0",
  2118 => x"00",
  2119 => x"7f",
  2120 => x"00",
  2121 => x"3e",
  2122 => x"61",
  2123 => x"00",
  2124 => x"fb",
  2125 => x"92",
  2126 => x"66",
  2127 => x"10",
  2128 => x"0c",
  2129 => x"28",
  2130 => x"00",
  2131 => x"55",
  2132 => x"01",
  2133 => x"fe",
  2134 => x"66",
  2135 => x"08",
  2136 => x"0c",
  2137 => x"28",
  2138 => x"00",
  2139 => x"aa",
  2140 => x"01",
  2141 => x"ff",
  2142 => x"67",
  2143 => x"0c",
  2144 => x"33",
  2145 => x"fc",
  2146 => x"f2",
  2147 => x"01",
  2148 => x"81",
  2149 => x"00",
  2150 => x"00",
  2151 => x"06",
  2152 => x"70",
  2153 => x"ff",
  2154 => x"4e",
  2155 => x"75",
  2156 => x"33",
  2157 => x"fc",
  2158 => x"02",
  2159 => x"04",
  2160 => x"81",
  2161 => x"00",
  2162 => x"00",
  2163 => x"06",
  2164 => x"0c",
  2165 => x"a8",
  2166 => x"46",
  2167 => x"41",
  2168 => x"54",
  2169 => x"31",
  2170 => x"00",
  2171 => x"36",
  2172 => x"66",
  2173 => x"24",
  2174 => x"13",
  2175 => x"fc",
  2176 => x"00",
  2177 => x"0c",
  2178 => x"00",
  2179 => x"7f",
  2180 => x"00",
  2181 => x"28",
  2182 => x"0c",
  2183 => x"a8",
  2184 => x"32",
  2185 => x"20",
  2186 => x"20",
  2187 => x"20",
  2188 => x"00",
  2189 => x"3a",
  2190 => x"67",
  2191 => x"36",
  2192 => x"13",
  2193 => x"fc",
  2194 => x"00",
  2195 => x"10",
  2196 => x"00",
  2197 => x"7f",
  2198 => x"00",
  2199 => x"28",
  2200 => x"0c",
  2201 => x"a8",
  2202 => x"36",
  2203 => x"20",
  2204 => x"20",
  2205 => x"20",
  2206 => x"00",
  2207 => x"3a",
  2208 => x"67",
  2209 => x"24",
  2210 => x"13",
  2211 => x"fc",
  2212 => x"00",
  2213 => x"00",
  2214 => x"00",
  2215 => x"7f",
  2216 => x"00",
  2217 => x"28",
  2218 => x"0c",
  2219 => x"a8",
  2220 => x"46",
  2221 => x"41",
  2222 => x"54",
  2223 => x"33",
  2224 => x"00",
  2225 => x"52",
  2226 => x"66",
  2227 => x"ac",
  2228 => x"0c",
  2229 => x"a8",
  2230 => x"32",
  2231 => x"20",
  2232 => x"20",
  2233 => x"20",
  2234 => x"00",
  2235 => x"56",
  2236 => x"66",
  2237 => x"a2",
  2238 => x"13",
  2239 => x"fc",
  2240 => x"00",
  2241 => x"20",
  2242 => x"00",
  2243 => x"7f",
  2244 => x"00",
  2245 => x"28",
  2246 => x"20",
  2247 => x"28",
  2248 => x"00",
  2249 => x"0a",
  2250 => x"c0",
  2251 => x"bc",
  2252 => x"00",
  2253 => x"ff",
  2254 => x"ff",
  2255 => x"00",
  2256 => x"0c",
  2257 => x"80",
  2258 => x"00",
  2259 => x"00",
  2260 => x"02",
  2261 => x"00",
  2262 => x"66",
  2263 => x"88",
  2264 => x"22",
  2265 => x"39",
  2266 => x"00",
  2267 => x"7f",
  2268 => x"00",
  2269 => x"3e",
  2270 => x"30",
  2271 => x"28",
  2272 => x"00",
  2273 => x"0e",
  2274 => x"e0",
  2275 => x"58",
  2276 => x"d2",
  2277 => x"80",
  2278 => x"23",
  2279 => x"c1",
  2280 => x"00",
  2281 => x"7f",
  2282 => x"00",
  2283 => x"42",
  2284 => x"0c",
  2285 => x"39",
  2286 => x"00",
  2287 => x"20",
  2288 => x"00",
  2289 => x"7f",
  2290 => x"00",
  2291 => x"28",
  2292 => x"66",
  2293 => x"24",
  2294 => x"20",
  2295 => x"28",
  2296 => x"00",
  2297 => x"2c",
  2298 => x"e0",
  2299 => x"58",
  2300 => x"48",
  2301 => x"40",
  2302 => x"e0",
  2303 => x"58",
  2304 => x"23",
  2305 => x"c0",
  2306 => x"00",
  2307 => x"7f",
  2308 => x"00",
  2309 => x"2a",
  2310 => x"20",
  2311 => x"28",
  2312 => x"00",
  2313 => x"24",
  2314 => x"e0",
  2315 => x"58",
  2316 => x"48",
  2317 => x"40",
  2318 => x"e0",
  2319 => x"58",
  2320 => x"d2",
  2321 => x"80",
  2322 => x"53",
  2323 => x"28",
  2324 => x"00",
  2325 => x"10",
  2326 => x"66",
  2327 => x"f8",
  2328 => x"60",
  2329 => x"32",
  2330 => x"70",
  2331 => x"00",
  2332 => x"23",
  2333 => x"c0",
  2334 => x"00",
  2335 => x"7f",
  2336 => x"00",
  2337 => x"2a",
  2338 => x"30",
  2339 => x"28",
  2340 => x"00",
  2341 => x"16",
  2342 => x"e0",
  2343 => x"58",
  2344 => x"d2",
  2345 => x"80",
  2346 => x"53",
  2347 => x"28",
  2348 => x"00",
  2349 => x"10",
  2350 => x"66",
  2351 => x"f8",
  2352 => x"23",
  2353 => x"c1",
  2354 => x"00",
  2355 => x"7f",
  2356 => x"00",
  2357 => x"2e",
  2358 => x"20",
  2359 => x"01",
  2360 => x"10",
  2361 => x"28",
  2362 => x"00",
  2363 => x"12",
  2364 => x"e1",
  2365 => x"48",
  2366 => x"10",
  2367 => x"28",
  2368 => x"00",
  2369 => x"11",
  2370 => x"33",
  2371 => x"c0",
  2372 => x"00",
  2373 => x"7f",
  2374 => x"00",
  2375 => x"4e",
  2376 => x"e8",
  2377 => x"48",
  2378 => x"d2",
  2379 => x"80",
  2380 => x"70",
  2381 => x"00",
  2382 => x"10",
  2383 => x"28",
  2384 => x"00",
  2385 => x"0d",
  2386 => x"33",
  2387 => x"c0",
  2388 => x"00",
  2389 => x"7f",
  2390 => x"00",
  2391 => x"4a",
  2392 => x"92",
  2393 => x"80",
  2394 => x"92",
  2395 => x"80",
  2396 => x"23",
  2397 => x"c1",
  2398 => x"00",
  2399 => x"7f",
  2400 => x"00",
  2401 => x"46",
  2402 => x"33",
  2403 => x"fc",
  2404 => x"02",
  2405 => x"05",
  2406 => x"81",
  2407 => x"00",
  2408 => x"00",
  2409 => x"06",
  2410 => x"70",
  2411 => x"00",
  2412 => x"4e",
  2413 => x"75",
  2414 => x"20",
  2415 => x"39",
  2416 => x"00",
  2417 => x"7f",
  2418 => x"00",
  2419 => x"2a",
  2420 => x"23",
  2421 => x"c0",
  2422 => x"00",
  2423 => x"7f",
  2424 => x"00",
  2425 => x"32",
  2426 => x"66",
  2427 => x"28",
  2428 => x"42",
  2429 => x"b9",
  2430 => x"00",
  2431 => x"7f",
  2432 => x"00",
  2433 => x"32",
  2434 => x"30",
  2435 => x"39",
  2436 => x"00",
  2437 => x"7f",
  2438 => x"00",
  2439 => x"4e",
  2440 => x"e8",
  2441 => x"48",
  2442 => x"33",
  2443 => x"c0",
  2444 => x"00",
  2445 => x"7f",
  2446 => x"00",
  2447 => x"36",
  2448 => x"20",
  2449 => x"39",
  2450 => x"00",
  2451 => x"7f",
  2452 => x"00",
  2453 => x"2e",
  2454 => x"23",
  2455 => x"c0",
  2456 => x"00",
  2457 => x"7f",
  2458 => x"00",
  2459 => x"38",
  2460 => x"4e",
  2461 => x"75",
  2462 => x"20",
  2463 => x"39",
  2464 => x"00",
  2465 => x"7f",
  2466 => x"00",
  2467 => x"32",
  2468 => x"32",
  2469 => x"39",
  2470 => x"00",
  2471 => x"7f",
  2472 => x"00",
  2473 => x"4a",
  2474 => x"33",
  2475 => x"c1",
  2476 => x"00",
  2477 => x"7f",
  2478 => x"00",
  2479 => x"36",
  2480 => x"e2",
  2481 => x"49",
  2482 => x"65",
  2483 => x"04",
  2484 => x"e3",
  2485 => x"88",
  2486 => x"60",
  2487 => x"f8",
  2488 => x"d0",
  2489 => x"b9",
  2490 => x"00",
  2491 => x"7f",
  2492 => x"00",
  2493 => x"46",
  2494 => x"23",
  2495 => x"c0",
  2496 => x"00",
  2497 => x"7f",
  2498 => x"00",
  2499 => x"38",
  2500 => x"4e",
  2501 => x"75",
  2502 => x"48",
  2503 => x"e7",
  2504 => x"20",
  2505 => x"20",
  2506 => x"24",
  2507 => x"49",
  2508 => x"61",
  2509 => x"00",
  2510 => x"fa",
  2511 => x"10",
  2512 => x"66",
  2513 => x"7a",
  2514 => x"74",
  2515 => x"0f",
  2516 => x"4a",
  2517 => x"10",
  2518 => x"67",
  2519 => x"74",
  2520 => x"70",
  2521 => x"0a",
  2522 => x"12",
  2523 => x"32",
  2524 => x"00",
  2525 => x"00",
  2526 => x"b2",
  2527 => x"30",
  2528 => x"00",
  2529 => x"00",
  2530 => x"67",
  2531 => x"0a",
  2532 => x"d2",
  2533 => x"3c",
  2534 => x"00",
  2535 => x"20",
  2536 => x"b2",
  2537 => x"30",
  2538 => x"00",
  2539 => x"00",
  2540 => x"66",
  2541 => x"36",
  2542 => x"51",
  2543 => x"c8",
  2544 => x"ff",
  2545 => x"ea",
  2546 => x"70",
  2547 => x"00",
  2548 => x"10",
  2549 => x"28",
  2550 => x"00",
  2551 => x"0b",
  2552 => x"33",
  2553 => x"c0",
  2554 => x"00",
  2555 => x"7f",
  2556 => x"00",
  2557 => x"3c",
  2558 => x"0c",
  2559 => x"39",
  2560 => x"00",
  2561 => x"20",
  2562 => x"00",
  2563 => x"7f",
  2564 => x"00",
  2565 => x"28",
  2566 => x"66",
  2567 => x"08",
  2568 => x"30",
  2569 => x"28",
  2570 => x"00",
  2571 => x"14",
  2572 => x"e0",
  2573 => x"58",
  2574 => x"48",
  2575 => x"40",
  2576 => x"30",
  2577 => x"28",
  2578 => x"00",
  2579 => x"1a",
  2580 => x"e0",
  2581 => x"58",
  2582 => x"23",
  2583 => x"c0",
  2584 => x"00",
  2585 => x"7f",
  2586 => x"00",
  2587 => x"32",
  2588 => x"4c",
  2589 => x"df",
  2590 => x"04",
  2591 => x"04",
  2592 => x"70",
  2593 => x"ff",
  2594 => x"4e",
  2595 => x"75",
  2596 => x"41",
  2597 => x"e8",
  2598 => x"00",
  2599 => x"20",
  2600 => x"51",
  2601 => x"ca",
  2602 => x"ff",
  2603 => x"aa",
  2604 => x"20",
  2605 => x"39",
  2606 => x"00",
  2607 => x"7f",
  2608 => x"00",
  2609 => x"38",
  2610 => x"52",
  2611 => x"80",
  2612 => x"23",
  2613 => x"c0",
  2614 => x"00",
  2615 => x"7f",
  2616 => x"00",
  2617 => x"38",
  2618 => x"53",
  2619 => x"79",
  2620 => x"00",
  2621 => x"7f",
  2622 => x"00",
  2623 => x"36",
  2624 => x"66",
  2625 => x"8a",
  2626 => x"61",
  2627 => x"10",
  2628 => x"67",
  2629 => x"06",
  2630 => x"61",
  2631 => x"00",
  2632 => x"ff",
  2633 => x"56",
  2634 => x"60",
  2635 => x"80",
  2636 => x"4c",
  2637 => x"df",
  2638 => x"04",
  2639 => x"04",
  2640 => x"70",
  2641 => x"00",
  2642 => x"4e",
  2643 => x"75",
  2644 => x"0c",
  2645 => x"39",
  2646 => x"00",
  2647 => x"20",
  2648 => x"00",
  2649 => x"7f",
  2650 => x"00",
  2651 => x"28",
  2652 => x"67",
  2653 => x"3e",
  2654 => x"0c",
  2655 => x"39",
  2656 => x"00",
  2657 => x"0c",
  2658 => x"00",
  2659 => x"7f",
  2660 => x"00",
  2661 => x"28",
  2662 => x"67",
  2663 => x"78",
  2664 => x"20",
  2665 => x"39",
  2666 => x"00",
  2667 => x"7f",
  2668 => x"00",
  2669 => x"32",
  2670 => x"e0",
  2671 => x"88",
  2672 => x"d0",
  2673 => x"b9",
  2674 => x"00",
  2675 => x"7f",
  2676 => x"00",
  2677 => x"42",
  2678 => x"61",
  2679 => x"00",
  2680 => x"f9",
  2681 => x"66",
  2682 => x"66",
  2683 => x"60",
  2684 => x"10",
  2685 => x"39",
  2686 => x"00",
  2687 => x"7f",
  2688 => x"00",
  2689 => x"35",
  2690 => x"d0",
  2691 => x"40",
  2692 => x"30",
  2693 => x"30",
  2694 => x"00",
  2695 => x"00",
  2696 => x"e0",
  2697 => x"58",
  2698 => x"23",
  2699 => x"c0",
  2700 => x"00",
  2701 => x"7f",
  2702 => x"00",
  2703 => x"32",
  2704 => x"80",
  2705 => x"bc",
  2706 => x"ff",
  2707 => x"ff",
  2708 => x"00",
  2709 => x"0f",
  2710 => x"b0",
  2711 => x"7c",
  2712 => x"ff",
  2713 => x"ff",
  2714 => x"4e",
  2715 => x"75",
  2716 => x"20",
  2717 => x"39",
  2718 => x"00",
  2719 => x"7f",
  2720 => x"00",
  2721 => x"32",
  2722 => x"ee",
  2723 => x"88",
  2724 => x"d0",
  2725 => x"b9",
  2726 => x"00",
  2727 => x"7f",
  2728 => x"00",
  2729 => x"42",
  2730 => x"61",
  2731 => x"00",
  2732 => x"f9",
  2733 => x"32",
  2734 => x"66",
  2735 => x"2c",
  2736 => x"10",
  2737 => x"39",
  2738 => x"00",
  2739 => x"7f",
  2740 => x"00",
  2741 => x"35",
  2742 => x"c0",
  2743 => x"7c",
  2744 => x"00",
  2745 => x"7f",
  2746 => x"d0",
  2747 => x"40",
  2748 => x"d0",
  2749 => x"40",
  2750 => x"20",
  2751 => x"30",
  2752 => x"00",
  2753 => x"00",
  2754 => x"e0",
  2755 => x"58",
  2756 => x"48",
  2757 => x"40",
  2758 => x"e0",
  2759 => x"58",
  2760 => x"23",
  2761 => x"c0",
  2762 => x"00",
  2763 => x"7f",
  2764 => x"00",
  2765 => x"32",
  2766 => x"80",
  2767 => x"bc",
  2768 => x"f0",
  2769 => x"00",
  2770 => x"00",
  2771 => x"07",
  2772 => x"b0",
  2773 => x"bc",
  2774 => x"ff",
  2775 => x"ff",
  2776 => x"ff",
  2777 => x"ff",
  2778 => x"4e",
  2779 => x"75",
  2780 => x"70",
  2781 => x"00",
  2782 => x"4e",
  2783 => x"75",
  2784 => x"2f",
  2785 => x"02",
  2786 => x"20",
  2787 => x"39",
  2788 => x"00",
  2789 => x"7f",
  2790 => x"00",
  2791 => x"32",
  2792 => x"22",
  2793 => x"00",
  2794 => x"d0",
  2795 => x"80",
  2796 => x"d0",
  2797 => x"81",
  2798 => x"22",
  2799 => x"00",
  2800 => x"e0",
  2801 => x"88",
  2802 => x"e4",
  2803 => x"88",
  2804 => x"d0",
  2805 => x"b9",
  2806 => x"00",
  2807 => x"7f",
  2808 => x"00",
  2809 => x"42",
  2810 => x"24",
  2811 => x"00",
  2812 => x"61",
  2813 => x"00",
  2814 => x"f8",
  2815 => x"e0",
  2816 => x"66",
  2817 => x"52",
  2818 => x"20",
  2819 => x"01",
  2820 => x"e2",
  2821 => x"88",
  2822 => x"c0",
  2823 => x"7c",
  2824 => x"01",
  2825 => x"ff",
  2826 => x"b0",
  2827 => x"7c",
  2828 => x"01",
  2829 => x"ff",
  2830 => x"66",
  2831 => x"14",
  2832 => x"10",
  2833 => x"30",
  2834 => x"00",
  2835 => x"00",
  2836 => x"c1",
  2837 => x"42",
  2838 => x"52",
  2839 => x"80",
  2840 => x"61",
  2841 => x"00",
  2842 => x"f8",
  2843 => x"c4",
  2844 => x"66",
  2845 => x"36",
  2846 => x"e1",
  2847 => x"4a",
  2848 => x"14",
  2849 => x"10",
  2850 => x"60",
  2851 => x"0a",
  2852 => x"14",
  2853 => x"30",
  2854 => x"00",
  2855 => x"00",
  2856 => x"e1",
  2857 => x"4a",
  2858 => x"14",
  2859 => x"30",
  2860 => x"00",
  2861 => x"01",
  2862 => x"e1",
  2863 => x"5a",
  2864 => x"c2",
  2865 => x"7c",
  2866 => x"00",
  2867 => x"01",
  2868 => x"67",
  2869 => x"02",
  2870 => x"e8",
  2871 => x"4a",
  2872 => x"c4",
  2873 => x"bc",
  2874 => x"00",
  2875 => x"00",
  2876 => x"0f",
  2877 => x"ff",
  2878 => x"23",
  2879 => x"c2",
  2880 => x"00",
  2881 => x"7f",
  2882 => x"00",
  2883 => x"32",
  2884 => x"84",
  2885 => x"bc",
  2886 => x"ff",
  2887 => x"ff",
  2888 => x"f0",
  2889 => x"0f",
  2890 => x"20",
  2891 => x"02",
  2892 => x"24",
  2893 => x"1f",
  2894 => x"b0",
  2895 => x"7c",
  2896 => x"ff",
  2897 => x"ff",
  2898 => x"4e",
  2899 => x"75",
  2900 => x"24",
  2901 => x"1f",
  2902 => x"70",
  2903 => x"00",
  2904 => x"4e",
  2905 => x"75",
  2906 => x"41",
  2907 => x"f9",
  2908 => x"00",
  2909 => x"7f",
  2910 => x"00",
  2911 => x"04",
  2912 => x"20",
  2913 => x"bc",
  2914 => x"12",
  2915 => x"34",
  2916 => x"56",
  2917 => x"78",
  2918 => x"21",
  2919 => x"7c",
  2920 => x"fe",
  2921 => x"dc",
  2922 => x"ba",
  2923 => x"98",
  2924 => x"00",
  2925 => x"04",
  2926 => x"21",
  2927 => x"7c",
  2928 => x"aa",
  2929 => x"55",
  2930 => x"cc",
  2931 => x"22",
  2932 => x"00",
  2933 => x"02",
  2934 => x"11",
  2935 => x"7c",
  2936 => x"00",
  2937 => x"33",
  2938 => x"00",
  2939 => x"03",
  2940 => x"11",
  2941 => x"7c",
  2942 => x"00",
  2943 => x"fe",
  2944 => x"00",
  2945 => x"04",
  2946 => x"20",
  2947 => x"10",
  2948 => x"22",
  2949 => x"28",
  2950 => x"00",
  2951 => x"04",
  2952 => x"90",
  2953 => x"bc",
  2954 => x"12",
  2955 => x"34",
  2956 => x"aa",
  2957 => x"33",
  2958 => x"92",
  2959 => x"bc",
  2960 => x"fe",
  2961 => x"22",
  2962 => x"ba",
  2963 => x"98",
  2964 => x"80",
  2965 => x"81",
  2966 => x"4e",
  2967 => x"75",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;

