
--
-- Copyright (c) 2008-2021 Sytse van Slooten
--
-- Permission is hereby granted to any person obtaining a copy of these VHDL source files and
-- other language source files and associated documentation files ("the materials") to use
-- these materials solely for personal, non-commercial purposes.
-- You are also granted permission to make changes to the materials, on the condition that this
-- copyright notice is retained unchanged.
--
-- The materials are distributed in the hope that they will be useful, but WITHOUT ANY WARRANTY;
-- without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
--

-- $Revision$

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity vgafont is
   port(
      ix : in std_logic_vector(15 downto 0);
      pix : out std_logic;
      vgaclk : in std_logic
   );
end vgafont;

architecture implementation of vgafont is

constant vga_font : std_logic_vector(0 to 32767) :=                          -- INSERT FONT HERE
   "0000000000000000100000000000000000000000000000000000000000000000"  &     -- 00000-00063 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 00064-00127 FONTDATA
   "0010000000000000100000000000000000000000000000000000000000000000"  &     -- 00128-00191 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 00192-00255 FONTDATA
   "0000000000000000100000000000000000000000000000000000000000000000"  &     -- 00256-00319 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 00320-00383 FONTDATA
   "0010000000010011100001110100000000000000000000000000000000000000"  &     -- 00384-00447 FONTDATA
   "0000000000000000000000000000001000000000000000000000000000000000"  &     -- 00448-00511 FONTDATA
   "0000000000010011100001110100000000000000000000000000000000000000"  &     -- 00512-00575 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 00576-00639 FONTDATA
   "0010000000000000100000000000000000000000000000000000000000000000"  &     -- 00640-00703 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 00704-00767 FONTDATA
   "0000000000000000100000000000000000000000000000000000000000000000"  &     -- 00768-00831 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 00832-00895 FONTDATA
   "0010000000000000100000000000000000000000000000000000000000000000"  &     -- 00896-00959 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 00960-01023 FONTDATA
   "0011101001100000100000000000000000000000000000000000000000000000"  &     -- 01024-01087 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 01088-01151 FONTDATA
   "0000110000000000100000000000000000000000000000000000000000000000"  &     -- 01152-01215 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 01216-01279 FONTDATA
   "0010110000000000100000000000000000100000000000000000000000000000"  &     -- 01280-01343 FONTDATA
   "0000000000000000000000000000001010000000000000000000000000000000"  &     -- 01344-01407 FONTDATA
   "0000110000010011100001110100000000001001000000000000000000000000"  &     -- 01408-01471 FONTDATA
   "0000000000000000000000000000001010000000000000000000000000000000"  &     -- 01472-01535 FONTDATA
   "0011110001110011100001110100000000000001000000000000000000000000"  &     -- 01536-01599 FONTDATA
   "0000000000000000000000000000001000000000000000000000000000000000"  &     -- 01600-01663 FONTDATA
   "0000000000000000100000000000000000100000000000000000000000000000"  &     -- 01664-01727 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 01728-01791 FONTDATA
   "0010000000000000100000000000000000000000000000000000000000000000"  &     -- 01792-01855 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 01856-01919 FONTDATA
   "0000000000000000100000000000000000000000000000000000000000000000"  &     -- 01920-01983 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 01984-02047 FONTDATA
   "0001111001100000000000000000000000000000000000000000010100000000"  &     -- 02048-02111 FONTDATA
   "0010111010011110101001111010000000100000100100000000000000000000"  &     -- 02112-02175 FONTDATA
   "0010000001000000000000000000000000000000000000001011010111000001"  &     -- 02176-02239 FONTDATA
   "1010111010011111111111111110001000100000100110000000000000000111"  &     -- 02240-02303 FONTDATA
   "0000000100000000000000000000001000100010010000001011011111000001"  &     -- 02304-02367 FONTDATA
   "1011111101011001111110000111011010100010100110000000000000000111"  &     -- 02368-02431 FONTDATA
   "0010000100010011000001110100001001001011010000001111011111000001"  &     -- 02432-02495 FONTDATA
   "1111111101101001111110000011010010001010010010000000100000001111"  &     -- 02496-02559 FONTDATA
   "0001000101110011000001110100001001000011100000001111111111000001"  &     -- 02560-02623 FONTDATA
   "1011111101100001111110000011011000001010010000000000000000011001"  &     -- 02624-02687 FONTDATA
   "0010000000000000000000000000000000100000100000001011110111000001"  &     -- 02688-02751 FONTDATA
   "1011011111110111111111111111011000001000001000000000000000010011"  &     -- 02752-02815 FONTDATA
   "0000000000000000000000000000000000000000000000000000010100000000"  &     -- 02816-02879 FONTDATA
   "0000011010110110000011111110000000000000001000000000000000010010"  &     -- 02880-02943 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 02944-03007 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 03008-03071 FONTDATA
   "0011111001000000000000000000000000000000000000001011010111000001"  &     -- 03072-03135 FONTDATA
   "1000000010000111010101111010001000000000000000000000000000000011"  &     -- 03136-03199 FONTDATA
   "0001100100100000000000000000001000011010000000001011011111000011"  &     -- 03200-03263 FONTDATA
   "1011111110011111111111111110001000100010100100000000000000000011"  &     -- 03264-03327 FONTDATA
   "0011100101000000000000000000001000111010000000000100001000000010"  &     -- 03328-03391 FONTDATA
   "0111111100011110101010000101000010100010100110000000100000000000"  &     -- 03392-03455 FONTDATA
   "0001000000110011000001110100000001001001110000000100100000000000"  &     -- 03456-03519 FONTDATA
   "0100000001000000000010000001000010000000010010000000100000011110"  &     -- 03520-03583 FONTDATA
   "0011000101010011000001110100001001011011110000000100100000000000"  &     -- 03584-03647 FONTDATA
   "0100100001100100000010000000010000001010010000000000000000011110"  &     -- 03648-03711 FONTDATA
   "0000000100000000000000000000011000111010000000001011100111001001"  &     -- 03712-03775 FONTDATA
   "1011111110110111111111111110011000001010001000000000000000000011"  &     -- 03776-03839 FONTDATA
   "0010000000000000000000000000010000000000000000001011000111001001"  &     -- 03840-03903 FONTDATA
   "1011011110010111111111111110001000000000001000000000000000000001"  &     -- 03904-03967 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 03968-04031 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 04032-04095 FONTDATA
   "0001111001000000010000000001000000001100000000001000011011000001"  &     -- 04096-04159 FONTDATA
   "1001000110000111010101110010000000000000000000000000000000000001"  &     -- 04160-04223 FONTDATA
   "0010000000100000010000000001001000011110000000001100011011000001"  &     -- 04224-04287 FONTDATA
   "1111111110011111111101111100000000100010100100000000000000000001"  &     -- 04288-04351 FONTDATA
   "0000000100000000010000000001001000110010100000000100100000000010"  &     -- 04352-04415 FONTDATA
   "0110111000011110101000001101000000100010100110000000100000000000"  &     -- 04416-04479 FONTDATA
   "0110000101110011010001110100000001001001100000000100100000110010"  &     -- 04480-04543 FONTDATA
   "0000000001000110000010000001000010000000000010000000100000011100"  &     -- 04544-04607 FONTDATA
   "0001000101010011010001110110010001010011010000000100100000111000"  &     -- 04608-04671 FONTDATA
   "0100000001100100000010001000010010001000000000000000000000011100"  &     -- 04672-04735 FONTDATA
   "0010000000000000010000000010010000111010010000001011100111001001"  &     -- 04736-04799 FONTDATA
   "1110100010110111111101111110010000001010000000000000000000000001"  &     -- 04800-04863 FONTDATA
   "0000000000000000010000000010000000001100000000001011000111000001"  &     -- 04864-04927 FONTDATA
   "1011111110010111111101110110000000000000000000000000000000000001"  &     -- 04928-04991 FONTDATA
   "0010000000000000010000000000000000000000000000000000000000000000"  &     -- 04992-05055 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 05056-05119 FONTDATA
   "0011101001000000010000000000110000011100000000001000011011000100"  &     -- 05120-05183 FONTDATA
   "1101000110000111010001110000100000000000000001101010110111100001"  &     -- 05184-05247 FONTDATA
   "0000011000000000010000000000011000011100001000001000111011000100"  &     -- 05248-05311 FONTDATA
   "1111111110011111111101111100100001110111100101111111111111100001"  &     -- 05312-05375 FONTDATA
   "0110011000100000010000000011011100010010101000000000100000000100"  &     -- 05376-05439 FONTDATA
   "0010111000011110101100001101000001111111110111010101101000100000"  &     -- 05440-05503 FONTDATA
   "0100011010010011010001110111010101011010100100000100000000111110"  &     -- 05504-05567 FONTDATA
   "0000000001000110000010001001000001111101010010111111100000111100"  &     -- 05568-05631 FONTDATA
   "0111011011010011010001110111010101010010010100000110100000111111"  &     -- 05632-05695 FONTDATA
   "0000011001110110000010001010010001111100111001111011110000111100"  &     -- 05696-05759 FONTDATA
   "0000000000000000010000000000010000010100011000011011100111000101"  &     -- 05760-05823 FONTDATA
   "1110100010110111111001111110010000011101101101111111111111100001"  &     -- 05824-05887 FONTDATA
   "0010000000000000010000000000010000010100001000011001000111000100"  &     -- 05888-05951 FONTDATA
   "1110100010000111111001110100000000000001001100000100001111100001"  &     -- 05952-06015 FONTDATA
   "0000000000000000010000000000000000000000000000000000000000000000"  &     -- 06016-06079 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 06080-06143 FONTDATA
   "0000000000000000000000000010101000001000000000001000111000000000"  &     -- 06144-06207 FONTDATA
   "1101000110000111010001110000000000010111000001010101010101100001"  &     -- 06208-06271 FONTDATA
   "0110000000000000000000000010101100011010000000001000111011000000"  &     -- 06272-06335 FONTDATA
   "1111111110011111111001110000100000111111100101111111011111110001"  &     -- 06336-06399 FONTDATA
   "0100000000000000000000000010101100010010101000000001011011001000"  &     -- 06400-06463 FONTDATA
   "0010111010011000101100001101100000101010100111101010101010010000"  &     -- 06464-06527 FONTDATA
   "0110000010010011000001110100111101001010101100001111011011001001"  &     -- 06528-06591 FONTDATA
   "0010011011010110101110001111000000000010110011000010100000011000"  &     -- 06592-06655 FONTDATA
   "0100000010010011000001110101111101010100011100010111111111000011"  &     -- 06656-06719 FONTDATA
   "1010011011110010101110001110010001101001010101000100010010101101"  &     -- 06720-06783 FONTDATA
   "0110000000000000000000000001100100010110011000011001111111000010"  &     -- 06784-06847 FONTDATA
   "1110100010100111111001110100010001111101101101111111011111100101"  &     -- 06848-06911 FONTDATA
   "0000000000000000000000000001100000000010000000001000000001000000"  &     -- 06912-06975 FONTDATA
   "1100100010000111010001110000000000010100101001111011001101000100"  &     -- 06976-07039 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 07040-07103 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 07104-07167 FONTDATA
   "0110000000000000000000000000000000000010001001001000101010000000"  &     -- 07168-07231 FONTDATA
   "1101000110000111010001110000000000011101000001010100010101000001"  &     -- 07232-07295 FONTDATA
   "0100000010000000000000000000101100011010001101001000101010001000"  &     -- 07296-07359 FONTDATA
   "1111111110011111111001110000000001111111100101111111011101000001"  &     -- 07360-07423 FONTDATA
   "0110000010000000000000000011111100011000101101000010100000001000"  &     -- 07424-07487 FONTDATA
   "0110111000011000101000001011100001100110100110101011101010000000"  &     -- 07488-07551 FONTDATA
   "0101111011110011000001110111010101001110101101011110100100000001"  &     -- 07552-07615 FONTDATA
   "1100000101010000000010011111100001000100010111000000100010110100"  &     -- 07616-07679 FONTDATA
   "0111111010110011000001110111100101011110011101010100100100000001"  &     -- 07680-07743 FONTDATA
   "1100011101110010001110001100010001001101010100000100010010110100"  &     -- 07744-07807 FONTDATA
   "0101111010100000000000000000100100011010011101001001111011000010"  &     -- 07808-07871 FONTDATA
   "1110100110100111011101110000010001101101101001111110011101000001"  &     -- 07872-07935 FONTDATA
   "0111111010100000000000000000100000000000001101001001111011000010"  &     -- 07936-07999 FONTDATA
   "1110100110000111010001110000000000100100101001111010001101000001"  &     -- 08000-08063 FONTDATA
   "0001101000100000000000000000000000000000001000000000000000000000"  &     -- 08064-08127 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 08128-08191 FONTDATA
   "0000000000000000000000000001010000000010000000001000001010000100"  &     -- 08192-08255 FONTDATA
   "1101000110100111010001110000000001011101000001010100010101000001"  &     -- 08256-08319 FONTDATA
   "0110000000000000000000000001111100010010000000001010001010000100"  &     -- 08320-08383 FONTDATA
   "1111111110111111111001111010000001111111100101111110011101000001"  &     -- 08384-08447 FONTDATA
   "0100000000000000000000000001111100010100101000010010000100001100"  &     -- 08448-08511 FONTDATA
   "0010111000011000101000001011000000100010100110101011101010100000"  &     -- 08512-08575 FONTDATA
   "0110111011010011000001110100010101001100101100010100000100001101"  &     -- 08576-08639 FONTDATA
   "1000000001000000000010011101100000000000010111000001100110111100"  &     -- 08640-08703 FONTDATA
   "0100000010010011000001110110110101010010011100000100100000000111"  &     -- 08704-08767 FONTDATA
   "1000000001110000000010001100110001001001010100000101010010011100"  &     -- 08768-08831 FONTDATA
   "0111000000100000000000000010110100011010011000001001111011000110"  &     -- 08832-08895 FONTDATA
   "1110100110110111011101111000010001101001101001111100011101000001"  &     -- 08896-08959 FONTDATA
   "0000000000000000000000000010010000001000000000001001011011000100"  &     -- 08960-09023 FONTDATA
   "1110100110000111011101110000000000100000101001111000001101000001"  &     -- 09024-09087 FONTDATA
   "0010010000000000000000000000000000000000000000000000000000000000"  &     -- 09088-09151 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 09152-09215 FONTDATA
   "0010000000011001001000111000000000010010000000001010001010000000"  &     -- 09216-09279 FONTDATA
   "1101000110100111010101010010000001011101000001010100010101000001"  &     -- 09280-09343 FONTDATA
   "0000000000011001001000111000111000010110001000011010001010000000"  &     -- 09344-09407 FONTDATA
   "1111111110111111111101111010000001111111100101111110011101100001"  &     -- 09408-09471 FONTDATA
   "0110000000011001001000111000111100010100101000010000000100000000"  &     -- 09472-09535 FONTDATA
   "0010111000011000101000111001000000100010100110101010101010100000"  &     -- 09536-09599 FONTDATA
   "0100111011011111001001111100000100011000100110000100000100111010"  &     -- 09600-09663 FONTDATA
   "0000000001000000010010010101000000000000010010000000100110011100"  &     -- 09664-09727 FONTDATA
   "0110111010011111001001111100100100010010010110000100100000111010"  &     -- 09728-09791 FONTDATA
   "1000000001100000000010111100110001001001010100000101010010011100"  &     -- 09792-09855 FONTDATA
   "0001111000100111001001011000100000011010011000001001111011000000"  &     -- 09856-09919 FONTDATA
   "1110100110110111011101111000110001101001101101111101011101000001"  &     -- 09920-09983 FONTDATA
   "0010010000000111001001011000000000011000001000001001011011000000"  &     -- 09984-10047 FONTDATA
   "0111110110010111011101010010000000100000101001111000001101000001"  &     -- 10048-10111 FONTDATA
   "0000010000000111001001011000000000000000000000000000000000000000"  &     -- 10112-10175 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 10176-10239 FONTDATA
   "0000000000011001001000111011010000001110000000011011011010000000"  &     -- 10240-10303 FONTDATA
   "1100000010100111010101011010000001011101000001010101010101100001"  &     -- 10304-10367 FONTDATA
   "0010000000011001001000111011111000011110000000011011011010000000"  &     -- 10368-10431 FONTDATA
   "1111111110111111111101011010000001111111100101111111010111100001"  &     -- 10432-10495 FONTDATA
   "0000000000011001001000111011101000010000000000000000000100000010"  &     -- 10496-10559 FONTDATA
   "0011111100011000101000110001000000100010100110101010101110000000"  &     -- 10560-10623 FONTDATA
   "0110111001011111001001111111001001001000110010100100000100110011"  &     -- 10624-10687 FONTDATA
   "0000000001000000010010100101000000000000010010000000101100011101"  &     -- 10688-10751 FONTDATA
   "0000000000011111001001111111100001010010110010100100100001111001"  &     -- 10752-10815 FONTDATA
   "0000100001100000010010110100010001001001010000000100011110011100"  &     -- 10816-10879 FONTDATA
   "0011000000100111001001011011100000011110000000001011111011001000"  &     -- 10880-10943 FONTDATA
   "0111110110111111011101011010110001111101101101111101111111100001"  &     -- 10944-11007 FONTDATA
   "0000010000000111001001011011000000001100000000001011011010000000"  &     -- 11008-11071 FONTDATA
   "0111010110011111011101011010100000110100101101111001100101100001"  &     -- 11072-11135 FONTDATA
   "0010000000000111001001011000000000000000000000000000000000000000"  &     -- 11136-11199 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 11200-11263 FONTDATA
   "0010000000000000000000000000001000000100000000000010000000000000"  &     -- 11264-11327 FONTDATA
   "0110111010011110101000001010000000000010100101000010000010100001"  &     -- 11328-11391 FONTDATA
   "0000000010000000000000000000101000011010000000001111011011000010"  &     -- 11392-11455 FONTDATA
   "1110111010111111111101011010000001111111100101111111010111100101"  &     -- 11456-11519 FONTDATA
   "0010000010000000000000000000101000011010010000001111011111010010"  &     -- 11520-11583 FONTDATA
   "1011111101111001111111010111010001111111110100111111010101100100"  &     -- 11584-11647 FONTDATA
   "0000111011001101000001101100001001001010010010101111111111010001"  &     -- 11648-11711 FONTDATA
   "1011111101101001110111100111010001111111010010011111111001101101"  &     -- 11712-11775 FONTDATA
   "0010000011001101000001101100101001011000100010101111111011000001"  &     -- 11776-11839 FONTDATA
   "1011110101101001010111010111010000110101010010011101101101111001"  &     -- 11840-11903 FONTDATA
   "0001000011100000000000000000101000011110100000001111111010001000"  &     -- 11904-11967 FONTDATA
   "1111010011011111011111011111010001111101111111111101110111110001"  &     -- 11968-12031 FONTDATA
   "0010000011000000000000000000000000000110000000000110100000001000"  &     -- 12032-12095 FONTDATA
   "0100010110011110001000001010000001001000101101100000010011110000"  &     -- 12096-12159 FONTDATA
   "0000010000000000000000000000000000000000000000000000000000000000"  &     -- 12160-12223 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 12224-12287 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 12288-12351 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000001"  &     -- 12352-12415 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 12416-12479 FONTDATA
   "0000000000000000000000000000000000000000001000001000000000000000"  &     -- 12480-12543 FONTDATA
   "0000000000000000000000000000000000000000000010000000000000000000"  &     -- 12544-12607 FONTDATA
   "0000000000000000000000000000000000000000001000001000000000000000"  &     -- 12608-12671 FONTDATA
   "0010000000001101000001101100000000001000000010000000000000000000"  &     -- 12672-12735 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000001000"  &     -- 12736-12799 FONTDATA
   "0000000000001101000001101100000000000000000000000000000000000000"  &     -- 12800-12863 FONTDATA
   "0000000000000000010000000000000000000001000000000100000000001000"  &     -- 12864-12927 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 12928-12991 FONTDATA
   "0000000000000000010000000000000000000001001000000100000001000000"  &     -- 12992-13055 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 13056-13119 FONTDATA
   "0000000000000000000000000000000000000000001000000000000001000000"  &     -- 13120-13183 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 13184-13247 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 13248-13311 FONTDATA
   "0010000000000000000100000000000000000000000000000000000000000000"  &     -- 13312-13375 FONTDATA
   "0000000000000000000000000000000000000001000000000000000000000000"  &     -- 13376-13439 FONTDATA
   "0000000000000000000100000000000000000000000000000000000000000000"  &     -- 13440-13503 FONTDATA
   "0000000000000000000000000000000000000001001000001000000000000000"  &     -- 13504-13567 FONTDATA
   "0010000000000000000100000000000000000000000000000000000000000000"  &     -- 13568-13631 FONTDATA
   "0000000000000000000000000000000000000000001000001000000000000000"  &     -- 13632-13695 FONTDATA
   "0000000000001101000101101100000000001000000000000000000000000000"  &     -- 13696-13759 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 13760-13823 FONTDATA
   "0010000000001101000101101100000000000000000000000000000000000000"  &     -- 13824-13887 FONTDATA
   "0000000000000000010000000000000000000001000000000100000000000000"  &     -- 13888-13951 FONTDATA
   "0000000000000000000100000000000000000000000000000000000000000000"  &     -- 13952-14015 FONTDATA
   "0000000000000000010000000000000000000001001000000100000001000000"  &     -- 14016-14079 FONTDATA
   "0010000000000000000100000000000000000000000000000000000000000000"  &     -- 14080-14143 FONTDATA
   "0000000000000000010000000000000000000000001000000000000001000000"  &     -- 14144-14207 FONTDATA
   "0000000000000000000100000000000000000000000000000000000000000000"  &     -- 14208-14271 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 14272-14335 FONTDATA
   "0000000000000000000100000000000000000000000000000000000000000000"  &     -- 14336-14399 FONTDATA
   "0000000000000000000000000000000100000000000000001000000001000000"  &     -- 14400-14463 FONTDATA
   "0010000000000000000100000000000000000000000000000000000000000000"  &     -- 14464-14527 FONTDATA
   "0000000000000000000000000000000100000001000000001000000001000000"  &     -- 14528-14591 FONTDATA
   "0000000000000000000100000000000000000000000000000000000000000000"  &     -- 14592-14655 FONTDATA
   "0000000000000000000000000000000100000001001000001000000001000000"  &     -- 14656-14719 FONTDATA
   "0010000000001101000101101100000000000000000000000000000000000000"  &     -- 14720-14783 FONTDATA
   "0000000000000000000000000000000100000001001000001100000001000000"  &     -- 14784-14847 FONTDATA
   "0000000000001101000101101100000000000000000000000000000000000000"  &     -- 14848-14911 FONTDATA
   "0000000000000000000000000000000100000001001000000100000001000000"  &     -- 14912-14975 FONTDATA
   "0010000000000000000100000000000000000000000000000000000000000000"  &     -- 14976-15039 FONTDATA
   "0000000000000000000000000000000100000000001000000100000000000000"  &     -- 15040-15103 FONTDATA
   "0000000000000000000100000000000000000000000000000000000000000000"  &     -- 15104-15167 FONTDATA
   "0000000000000000000000000000000100000000000000000100000000000000"  &     -- 15168-15231 FONTDATA
   "0010000000000000000100000000000000000000000000000000000000000000"  &     -- 15232-15295 FONTDATA
   "0000000000000000000000000000000100000000000000000000000000000000"  &     -- 15296-15359 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 15360-15423 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 15424-15487 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 15488-15551 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 15552-15615 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 15616-15679 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 15680-15743 FONTDATA
   "0000000000001101000001101100000000000000000000000000000000000000"  &     -- 15744-15807 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 15808-15871 FONTDATA
   "0010000000001101000001101100000000000000000000000000000000000000"  &     -- 15872-15935 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 15936-15999 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16000-16063 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16064-16127 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 16128-16191 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16192-16255 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16256-16319 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16320-16383 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16384-16447 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16448-16511 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 16512-16575 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16576-16639 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16640-16703 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16704-16767 FONTDATA
   "0010000000001101000001101100000000000000000000000000000000000000"  &     -- 16768-16831 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16832-16895 FONTDATA
   "0000000000001101000001101100000000000000000000000000000000000000"  &     -- 16896-16959 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 16960-17023 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 17024-17087 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 17088-17151 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 17152-17215 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 17216-17279 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 17280-17343 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 17344-17407 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 17408-17471 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 17472-17535 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 17536-17599 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 17600-17663 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 17664-17727 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 17728-17791 FONTDATA
   "0000000000001101000001101100000000000000000000000000000000000000"  &     -- 17792-17855 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 17856-17919 FONTDATA
   "0010000000001101000001101100000000000000000000000000000000000000"  &     -- 17920-17983 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 17984-18047 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 18048-18111 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 18112-18175 FONTDATA
   "0010000000000000000000000000000000000000000000000000000000000000"  &     -- 18176-18239 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 18240-18303 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 18304-18367 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 18368-18431 FONTDATA
   "0000000000000000000010000000000000000000000000000000000000000000"  &     -- 18432-18495 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 18496-18559 FONTDATA
   "0010000000000000000010000000000000000000000000000000000000000000"  &     -- 18560-18623 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 18624-18687 FONTDATA
   "0000000000000000000010000000000000000000000000000000000000000000"  &     -- 18688-18751 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 18752-18815 FONTDATA
   "0010000000001101000011101100000000000000000000000000000000000000"  &     -- 18816-18879 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 18880-18943 FONTDATA
   "0000000000001101000011101100000000000000000000000000000000000000"  &     -- 18944-19007 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 19008-19071 FONTDATA
   "0010000000000000000010000000000000000000000000000000000000000000"  &     -- 19072-19135 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 19136-19199 FONTDATA
   "0000000000000000000010000000000000000000000000000000000000000000"  &     -- 19200-19263 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 19264-19327 FONTDATA
   "0010000000000000000010000000000000000000000000000000000000000000"  &     -- 19328-19391 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 19392-19455 FONTDATA
   "0010000000000000000010000000000000000000000000000000000000000000"  &     -- 19456-19519 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 19520-19583 FONTDATA
   "0000000000000000000010000000000000000000000000000000000000000000"  &     -- 19584-19647 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 19648-19711 FONTDATA
   "0010000000000000000010000000000000000000000000000000000000000000"  &     -- 19712-19775 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 19776-19839 FONTDATA
   "0000000000001101000011101100000000000000000000000000000000000000"  &     -- 19840-19903 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 19904-19967 FONTDATA
   "0010000000001101000011101100000000000000000000000000000000000000"  &     -- 19968-20031 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20032-20095 FONTDATA
   "0000000000000000000010000000000000000000000000000000000000000000"  &     -- 20096-20159 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20160-20223 FONTDATA
   "0010000000000000000010000000000000000000000000000000000000000000"  &     -- 20224-20287 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20288-20351 FONTDATA
   "0000000000000000000010000000000000000000000000000000000000000000"  &     -- 20352-20415 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20416-20479 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20480-20543 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20544-20607 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20608-20671 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20672-20735 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20736-20799 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20800-20863 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20864-20927 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20928-20991 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 20992-21055 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21056-21119 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21120-21183 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21184-21247 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21248-21311 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21312-21375 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21376-21439 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21440-21503 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21504-21567 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21568-21631 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21632-21695 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21696-21759 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21760-21823 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21824-21887 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21888-21951 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 21952-22015 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22016-22079 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22080-22143 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22144-22207 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22208-22271 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22272-22335 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22336-22399 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22400-22463 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22464-22527 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22528-22591 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22592-22655 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22656-22719 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22720-22783 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22784-22847 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22848-22911 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22912-22975 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 22976-23039 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23040-23103 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23104-23167 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23168-23231 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23232-23295 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23296-23359 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23360-23423 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23424-23487 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23488-23551 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23552-23615 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23616-23679 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23680-23743 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23744-23807 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23808-23871 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23872-23935 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 23936-23999 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24000-24063 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24064-24127 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24128-24191 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24192-24255 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24256-24319 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24320-24383 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24384-24447 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24448-24511 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24512-24575 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24576-24639 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24640-24703 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24704-24767 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24768-24831 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24832-24895 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24896-24959 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 24960-25023 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25024-25087 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25088-25151 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25152-25215 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25216-25279 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25280-25343 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25344-25407 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25408-25471 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25472-25535 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25536-25599 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25600-25663 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25664-25727 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25728-25791 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25792-25855 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25856-25919 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25920-25983 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 25984-26047 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26048-26111 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26112-26175 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26176-26239 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26240-26303 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26304-26367 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26368-26431 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26432-26495 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26496-26559 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26560-26623 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26624-26687 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26688-26751 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26752-26815 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26816-26879 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26880-26943 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 26944-27007 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27008-27071 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27072-27135 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27136-27199 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27200-27263 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27264-27327 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27328-27391 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27392-27455 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27456-27519 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27520-27583 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27584-27647 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27648-27711 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27712-27775 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27776-27839 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27840-27903 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27904-27967 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 27968-28031 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28032-28095 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28096-28159 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28160-28223 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28224-28287 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28288-28351 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28352-28415 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28416-28479 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28480-28543 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28544-28607 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28608-28671 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28672-28735 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28736-28799 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28800-28863 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28864-28927 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28928-28991 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 28992-29055 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29056-29119 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29120-29183 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29184-29247 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29248-29311 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29312-29375 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29376-29439 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29440-29503 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29504-29567 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29568-29631 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29632-29695 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29696-29759 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29760-29823 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29824-29887 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29888-29951 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 29952-30015 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30016-30079 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30080-30143 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30144-30207 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30208-30271 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30272-30335 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30336-30399 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30400-30463 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30464-30527 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30528-30591 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30592-30655 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30656-30719 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30720-30783 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30784-30847 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30848-30911 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30912-30975 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 30976-31039 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31040-31103 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31104-31167 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31168-31231 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31232-31295 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31296-31359 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31360-31423 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31424-31487 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31488-31551 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31552-31615 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31616-31679 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31680-31743 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31744-31807 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31808-31871 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31872-31935 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 31936-31999 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32000-32063 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32064-32127 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32128-32191 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32192-32255 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32256-32319 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32320-32383 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32384-32447 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32448-32511 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32512-32575 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32576-32639 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"  &     -- 32640-32703 FONTDATA
   "0000000000000000000000000000000000000000000000000000000000000000"        -- 32704-32767 FONTDATA
;


begin
   process(vgaclk)
   begin
      if vgaclk='1' and vgaclk'event then
         pix <= vga_font(conv_integer(ix));
      end if;
   end process;
end implementation;

