--===========================================================================--
--
--  S Y N T H E Z I A B L E    SWTBUG ROM   C O R E
--
--  www.OpenCores.Org - April 2003
--  This core adheres to the GNU public license  
--
-- File name      : cfboot00.vhd
--
-- entity name    : boot_rom
--
-- Purpose        : Implements a 256 x 8 ROM containing the
--                  a boot program for Compact Flash
--                  SWTBUG is assumed to reside at
--                  LBA Address $F478 - $F479 of the Compact Flash
--                  Compact Flash is mapped at $8010
--                  ROM Map Switch at $8030 (clear for RAM)
--                  The idea of using a compact flash Boot ROM
--                  Is to save space in the FPGA rather by booting
--                  the ROM into RAM.
--                  
-- Dependencies   : ieee.Std_Logic_1164
--                  ieee.std_logic_unsigned
--                  ieee.std_logic_arith
--
-- Author         : John E. Kent      
--
--===========================================================================----
--
-- Revision History:
--
-- Date:          Revision         Author
-- 11 Apr 2003    0.1              John Kent
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity boot_rom is
  port (
    addr   : in   std_logic_vector(7 downto 0);
    data   : out  std_logic_vector(7 downto 0)
  );
end entity boot_rom;

architecture basic of boot_rom is
  constant width   : integer := 8;
  constant memsize : integer := 256;

  type rom_array is array(0 to memsize-1) of std_logic_vector(width-1 downto 0);

  constant rom_data : rom_array :=
(
"10001110", -- LDS #$A7FE
"10100111",
"11111110",
------------------
"11001110", -- LDX #$FF23
"11111111",
"00100011",
------------------
-- "11001110", -- LDX #$DF23
-- "11011111",
-- "00100011",
------------------
"11011111", -- STX $0004
"00000100",
"11001110", -- LDX #$1000
"00010000",
"00000000",
"11011111", -- STX $0006
"00000110",
"11000110", -- LDAB #$C0
"11000000",
"11011110", -- LDX $0004 *** MOVELP
"00000100",
"10100110", -- LDAA 0,X
"00000000",
"00001000", -- INX
"11011111", -- STX $0004
"00000100",
"11011110", -- LDX $0006
"00000110",
"10100111", -- STAA 0,X
"00000000",
"00001000", -- INX
"11011111", -- STX $0006
"00000110",
"01011010", -- DECB
"00100110", -- BNE MOVELP
"11101111",
"01111110", -- JMP $1000
"00010000",
"00000000",
--------------
"11001110", -- LDX #$E000
"11100000",
"00000000",
--------------
-- "11001110", -- LDX #$C000
-- "11000000",
-- "00000000",
--------------
"11011111", -- STX $0000
"00000000",
"11000110", -- LDAB #$78
"01111000",
"11010111", -- STAB $0003
"00000011",
"11001110", -- LDX #$8010
"10000000",
"00010000",
"10001101", -- BSR WAITRDY
"01011001",
"10000110", -- LDAA #$E0  (SELECT LBA MODE)
"11100000",
"10100111", -- STAA 6,X
"00000110",
"10001101", -- BSR WAITRDY
"01010011",
"10000110", -- LDAA #$01 (8 BIT I/O MODE)
"00000001",
"10100111", -- STAA 1,X
"00000001",
"10000110", -- LDAA #$EF (SET CONFIG COMMAND)
"11101111",
"10100111", -- STAA 7,X  (COMMAND REGISTER)
"00000111",
"11001110", -- LDX #$8010 *** RDLP1
"10000000",
"00010000",
"10001101", -- BSR WAITRDY
"01000110",
"10000110", -- LDAA #$01
"00000001",
"10100111", -- STAA 2,X (SECTOR COUNT)
"00000010",
"10010110", -- LDAA $0003
"00000011",
"10100111", -- STAA 3,X (SECTOR NUMBER)
"00000011",
"10000110", -- LDAA #$F4
"11110100",
"10100111", -- STAA 4,X (CYLINDER LOW)
"00000100",
"10000110", -- LDAA #$00
"00000000",
"10100111", -- STAA 5,X (CYLINDER HI)
"00000101",
"10000110", -- LDAA #$20 (READ SECTOR COMMAND)
"00100000",
"10100111", -- STAA 7,X (COMMAND REGISTER)
"00000111",
"10001101", -- BSR WAITRDY
"00110000",
"11000110", -- LDAB #$02
"00000010",
"11010111", -- STAB $0002 (HI BYTE COUNTER)
"00000010",
"01011111", -- CLRB
"11001110", -- LDX #$8010 *** RDLP2
"10000000",
"00010000",
"10100110", -- LDAA 7,X (STATUS REGISTER) *** WAITDRQ
"00000111",
"10000101", -- BITA #$08
"00001000",
"00100111", -- BEQ WAITDRQ
"11111010",
"10100110", -- LDAA 0,X (DATA REGISTER)
"00000000",
"11011110", -- LDX $0000 (LOAD ADDRESS)
"00000000",
"10100111", -- STAA 0,X
"00000000",
"00001000", -- INX
"11011111", -- STX $0000
"00000000",
"01011010", -- DECB
"00100110", -- BNE RDLP2
"11101011",
"01111010", -- DEC $0002 (HI BYTE COUNT)
"00000000",
"00000010",
"00100110", -- BNE RDLP2
"11100110",
"11010110", -- LDAB $0003 (LO SECTOR NUMBER)
"00000011",
"01011100", -- INCB
"11010111", -- STAB $0003
"00000011",
"11000001", -- CMPB #$7A
"01111010",
"00100110", -- BNE RDLP1
"10111101",
---------------------------------
-- "01111111", -- CLR $8030 (MAP SWITCH)
-- "10000000",
-- "00110000",
-- "11111110", -- LDX $FFFE
-- "11111111",
-- "11111110",
-- "01101110", -- JMP 0,X
-- "00000000",
--------------------------------
"00100000", -- BRA MOVE2
"00010001",
"00000001", -- NOP
"00000001", -- NOP
"00000001", -- NOP
"00000001", -- NOP
"00000001", -- NOP
"00000001", -- NOP
--------------------------------
"10100110", -- LDAA 7,X (STATUS REG) *** WAITRDY
"00000111",
"00101011", -- BMI WAITDRDY (BUSY = B7)
"11111100",
"10100110", -- LDAA 7,X
"00000111",
"10000101", -- BITA #$40
"01000000",
"00100111", -- BEQ WAITRDY
"11110110",
"00111001", -- RTS
--------------------------------
"11001110", -- LDX #$E3F8 *** MOVE2
"11100011",
"11111000",
"11011111", -- STX $0004
"00000100",
"11001110", -- LDX #$FFF8
"11111111",
"11111000",
"11011111", -- STX $0006
"00000110",
"11000110", -- LDAB #$08
"01110010",
"11011110", -- LDX $0004 *** MOVELP
"00000100",
"10100110", -- LDAA 0,X
"00000000",
"00001000", -- INX
"11011111", -- STX $0004
"00000100",
"11011110", -- LDX $0006
"00000110",
"10100111", -- STAA 0,X
"00000000",
"00001000", -- INX
"11011111", -- STX $0006
"00000110",
"01011010", -- DECB
"00100110", -- BNE MOVELP
"11101111",
"01111111", -- CLR $8030 (MAP SWITCH)
"10000000",
"00110000",
"11111110", -- LDX $FFFE
"11111111",
"11111110",
"01101110", -- JMP 0,X
"00000000",
--------------------------
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000",
"11111111",
"00000000"
);
begin
   data <= rom_data(conv_integer(addr)); 
end architecture basic;

