//
module char_rom(addr, data);
   
   input [9:0] addr;
   output reg [7:0] data;

   always @(addr)
     case (addr)

       	// char 0, '.'
	0: data <= 8'h00;
	1: data <= 8'h00;
	2: data <= 8'h00;
	3: data <= 8'h00;
	4: data <= 8'h00;
	5: data <= 8'h00;
	6: data <= 8'h00;
	7: data <= 8'h00;
	// char 1, '.'
	8: data <= 8'h00;
	9: data <= 8'h00;
	10: data <= 8'h00;
	11: data <= 8'h00;
	12: data <= 8'h00;
	13: data <= 8'h00;
	14: data <= 8'h00;
	15: data <= 8'h00;
	// char 2, '.'
	16: data <= 8'h00;
	17: data <= 8'h00;
	18: data <= 8'h00;
	19: data <= 8'h00;
	20: data <= 8'h00;
	21: data <= 8'h00;
	22: data <= 8'h00;
	23: data <= 8'h00;
	// char 3, '.'
	24: data <= 8'h00;
	25: data <= 8'h00;
	26: data <= 8'h00;
	27: data <= 8'h00;
	28: data <= 8'h00;
	29: data <= 8'h00;
	30: data <= 8'h00;
	31: data <= 8'h00;
	// char 4, '.'
	32: data <= 8'h00;
	33: data <= 8'h00;
	34: data <= 8'h00;
	35: data <= 8'h00;
	36: data <= 8'h00;
	37: data <= 8'h00;
	38: data <= 8'h00;
	39: data <= 8'h00;
	// char 5, '.'
	40: data <= 8'h00;
	41: data <= 8'h00;
	42: data <= 8'h00;
	43: data <= 8'h00;
	44: data <= 8'h00;
	45: data <= 8'h00;
	46: data <= 8'h00;
	47: data <= 8'h00;
	// char 6, '.'
	48: data <= 8'h00;
	49: data <= 8'h00;
	50: data <= 8'h00;
	51: data <= 8'h00;
	52: data <= 8'h00;
	53: data <= 8'h00;
	54: data <= 8'h00;
	55: data <= 8'h00;
	// char 7, '.'
	56: data <= 8'h00;
	57: data <= 8'h00;
	58: data <= 8'h00;
	59: data <= 8'h00;
	60: data <= 8'h00;
	61: data <= 8'h00;
	62: data <= 8'h00;
	63: data <= 8'h00;
	// char 8, '.'
	64: data <= 8'h00;
	65: data <= 8'h00;
	66: data <= 8'h00;
	67: data <= 8'h00;
	68: data <= 8'h00;
	69: data <= 8'h00;
	70: data <= 8'h00;
	71: data <= 8'h00;
	// char 9, '.'
	72: data <= 8'h00;
	73: data <= 8'h00;
	74: data <= 8'h00;
	75: data <= 8'h00;
	76: data <= 8'h00;
	77: data <= 8'h00;
	78: data <= 8'h00;
	79: data <= 8'h00;
	// char 10, '.'
	80: data <= 8'h00;
	81: data <= 8'h00;
	82: data <= 8'h00;
	83: data <= 8'h00;
	84: data <= 8'h00;
	85: data <= 8'h00;
	86: data <= 8'h00;
	87: data <= 8'h00;
	// char 11, '.'
	88: data <= 8'h00;
	89: data <= 8'h00;
	90: data <= 8'h00;
	91: data <= 8'h00;
	92: data <= 8'h00;
	93: data <= 8'h00;
	94: data <= 8'h00;
	95: data <= 8'h00;
	// char 12, '.'
	96: data <= 8'h00;
	97: data <= 8'h00;
	98: data <= 8'h00;
	99: data <= 8'h00;
	100: data <= 8'h00;
	101: data <= 8'h00;
	102: data <= 8'h00;
	103: data <= 8'h00;
	// char 13, '.'
	104: data <= 8'h00;
	105: data <= 8'h00;
	106: data <= 8'h00;
	107: data <= 8'h00;
	108: data <= 8'h00;
	109: data <= 8'h00;
	110: data <= 8'h00;
	111: data <= 8'h00;
	// char 14, '.'
	112: data <= 8'h00;
	113: data <= 8'h00;
	114: data <= 8'h00;
	115: data <= 8'h00;
	116: data <= 8'h00;
	117: data <= 8'h00;
	118: data <= 8'h00;
	119: data <= 8'h00;
	// char 15, '.'
	120: data <= 8'h00;
	121: data <= 8'h00;
	122: data <= 8'h00;
	123: data <= 8'h00;
	124: data <= 8'h00;
	125: data <= 8'h00;
	126: data <= 8'h00;
	127: data <= 8'h00;
	// char 16, '.'
	128: data <= 8'h00;
	129: data <= 8'h00;
	130: data <= 8'h00;
	131: data <= 8'h00;
	132: data <= 8'h00;
	133: data <= 8'h00;
	134: data <= 8'h00;
	135: data <= 8'h00;
	// char 17, '.'
	136: data <= 8'h00;
	137: data <= 8'h00;
	138: data <= 8'h00;
	139: data <= 8'h00;
	140: data <= 8'h00;
	141: data <= 8'h00;
	142: data <= 8'h00;
	143: data <= 8'h00;
	// char 18, '.'
	144: data <= 8'h00;
	145: data <= 8'h00;
	146: data <= 8'h00;
	147: data <= 8'h00;
	148: data <= 8'h00;
	149: data <= 8'h00;
	150: data <= 8'h00;
	151: data <= 8'h00;
	// char 19, '.'
	152: data <= 8'h00;
	153: data <= 8'h00;
	154: data <= 8'h00;
	155: data <= 8'h00;
	156: data <= 8'h00;
	157: data <= 8'h00;
	158: data <= 8'h00;
	159: data <= 8'h00;
	// char 20, '.'
	160: data <= 8'h00;
	161: data <= 8'h00;
	162: data <= 8'h00;
	163: data <= 8'h00;
	164: data <= 8'h00;
	165: data <= 8'h00;
	166: data <= 8'h00;
	167: data <= 8'h00;
	// char 21, '.'
	168: data <= 8'h00;
	169: data <= 8'h00;
	170: data <= 8'h00;
	171: data <= 8'h00;
	172: data <= 8'h00;
	173: data <= 8'h00;
	174: data <= 8'h00;
	175: data <= 8'h00;
	// char 22, '.'
	176: data <= 8'h00;
	177: data <= 8'h00;
	178: data <= 8'h00;
	179: data <= 8'h00;
	180: data <= 8'h00;
	181: data <= 8'h00;
	182: data <= 8'h00;
	183: data <= 8'h00;
	// char 23, '.'
	184: data <= 8'h00;
	185: data <= 8'h00;
	186: data <= 8'h00;
	187: data <= 8'h00;
	188: data <= 8'h00;
	189: data <= 8'h00;
	190: data <= 8'h00;
	191: data <= 8'h00;
	// char 24, '.'
	192: data <= 8'h00;
	193: data <= 8'h00;
	194: data <= 8'h00;
	195: data <= 8'h00;
	196: data <= 8'h00;
	197: data <= 8'h00;
	198: data <= 8'h00;
	199: data <= 8'h00;
	// char 25, '.'
	200: data <= 8'h00;
	201: data <= 8'h00;
	202: data <= 8'h00;
	203: data <= 8'h00;
	204: data <= 8'h00;
	205: data <= 8'h00;
	206: data <= 8'h00;
	207: data <= 8'h00;
	// char 26, '.'
	208: data <= 8'h00;
	209: data <= 8'h00;
	210: data <= 8'h00;
	211: data <= 8'h00;
	212: data <= 8'h00;
	213: data <= 8'h00;
	214: data <= 8'h00;
	215: data <= 8'h00;
	// char 27, '.'
	216: data <= 8'h00;
	217: data <= 8'h00;
	218: data <= 8'h00;
	219: data <= 8'h00;
	220: data <= 8'h00;
	221: data <= 8'h00;
	222: data <= 8'h00;
	223: data <= 8'h00;
	// char 28, '.'
	224: data <= 8'h00;
	225: data <= 8'h00;
	226: data <= 8'h00;
	227: data <= 8'h00;
	228: data <= 8'h00;
	229: data <= 8'h00;
	230: data <= 8'h00;
	231: data <= 8'h00;
	// char 29, '.'
	232: data <= 8'h00;
	233: data <= 8'h00;
	234: data <= 8'h00;
	235: data <= 8'h00;
	236: data <= 8'h00;
	237: data <= 8'h00;
	238: data <= 8'h00;
	239: data <= 8'h00;
	// char 30, '.'
	240: data <= 8'h00;
	241: data <= 8'h00;
	242: data <= 8'h00;
	243: data <= 8'h00;
	244: data <= 8'h00;
	245: data <= 8'h00;
	246: data <= 8'h00;
	247: data <= 8'h00;
	// char 31, '.'
	248: data <= 8'h00;
	249: data <= 8'h00;
	250: data <= 8'h00;
	251: data <= 8'h00;
	252: data <= 8'h00;
	253: data <= 8'h00;
	254: data <= 8'h00;
	255: data <= 8'h00;
	// char 32, ' '
	256: data <= 8'h00;
	257: data <= 8'h00;
	258: data <= 8'h00;
	259: data <= 8'h00;
	260: data <= 8'h00;
	261: data <= 8'h00;
	262: data <= 8'h00;
	263: data <= 8'h00;
	// char 33, '!'
	264: data <= 8'h10;
	265: data <= 8'h38;
	266: data <= 8'h38;
	267: data <= 8'h10;
	268: data <= 8'h10;
	269: data <= 8'h00;
	270: data <= 8'h10;
	271: data <= 8'h00;
	// char 34, '"'
	272: data <= 8'h6c;
	273: data <= 8'h6c;
	274: data <= 8'h48;
	275: data <= 8'h00;
	276: data <= 8'h00;
	277: data <= 8'h00;
	278: data <= 8'h00;
	279: data <= 8'h00;
	// char 35, '#'
	280: data <= 8'h00;
	281: data <= 8'h28;
	282: data <= 8'h7c;
	283: data <= 8'h28;
	284: data <= 8'h28;
	285: data <= 8'h7c;
	286: data <= 8'h28;
	287: data <= 8'h00;
	// char 36, '$'
	288: data <= 8'h10;  // ...X.... 10
	289: data <= 8'h7e;  // .XXXXXX. 7e
	290: data <= 8'h90;  // X..X.... 90
	291: data <= 8'h7c;  // .XXXXX.. 7c
	292: data <= 8'h12;  // ...X..X. 12
	293: data <= 8'hfc;  // XXXXXX.. fc
	294: data <= 8'h10;  // ...X.... 10
	295: data <= 8'h00;  // ........ 00
	// char 37, '%'
	296: data <= 8'h62;  // .XX...X. 62
	297: data <= 8'h94;  // X..X.X.. 94
	298: data <= 8'h68;  // .XX.X... 68
	299: data <= 8'h10;  // ...X.... 10
	300: data <= 8'h26;  // ..X..XX. 26
	301: data <= 8'h49;  // .X..X..X 49
	302: data <= 8'h86;  // X....XX. 86
	303: data <= 8'h00;  // ........ 00
	// char 38, '&'
	304: data <= 8'h30;  // ..XX.... 30
	305: data <= 8'h48;  // .X..X... 48
	306: data <= 8'h30;  // ..XX.... 30
	307: data <= 8'h48;  // .X..X... 48
	308: data <= 8'h85;  // X....X.X 85
	309: data <= 8'h46;  // .X...XX. 46
	310: data <= 8'h39;  // ..XXX..X 39
	311: data <= 8'h00;  // ........ 00
	// char 39, '''
	312: data <= 8'h30;
	313: data <= 8'h30;
	314: data <= 8'h20;
	315: data <= 8'h00;
	316: data <= 8'h00;
	317: data <= 8'h00;
	318: data <= 8'h00;
	319: data <= 8'h00;
	// char 40, '('
	320: data <= 8'h10;
	321: data <= 8'h20;
	322: data <= 8'h20;
	323: data <= 8'h20;
	324: data <= 8'h20;
	325: data <= 8'h20;
	326: data <= 8'h10;
	327: data <= 8'h00;
	// char 41, ')'
	328: data <= 8'h20;
	329: data <= 8'h10;
	330: data <= 8'h10;
	331: data <= 8'h10;
	332: data <= 8'h10;
	333: data <= 8'h10;
	334: data <= 8'h20;
	335: data <= 8'h00;
	// char 42, '*'
	336: data <= 8'h99;  // X..XX..X 00
	337: data <= 8'h5a;  // .X.XX.X. 00
	338: data <= 8'h3c;  // ..XXXX.. 00
	339: data <= 8'hff;  // XXXXXXXX 00
	340: data <= 8'h3c;  // ..XXXX.. 00
	341: data <= 8'h5a;  // .X.XX.X. 00
	342: data <= 8'h99;  // X..XX..X 00
	343: data <= 8'h00;  // ........ 00
	// char 43, '+'
	344: data <= 8'h00;
	345: data <= 8'h10;
	346: data <= 8'h10;
	347: data <= 8'h7c;
	348: data <= 8'h10;
	349: data <= 8'h10;
	350: data <= 8'h00;
	351: data <= 8'h00;
	// char 44, ','
	352: data <= 8'h00;
	353: data <= 8'h00;
	354: data <= 8'h00;
	355: data <= 8'h00;
	356: data <= 8'h00;
	357: data <= 8'h30;
	358: data <= 8'h30;
	359: data <= 8'h20;
	// char 45, '-'
	360: data <= 8'h00;
	361: data <= 8'h00;
	362: data <= 8'h00;
	363: data <= 8'h7c;
	364: data <= 8'h00;
	365: data <= 8'h00;
	366: data <= 8'h00;
	367: data <= 8'h00;
	// char 46, '.'
	368: data <= 8'h00;
	369: data <= 8'h00;
	370: data <= 8'h00;
	371: data <= 8'h00;
	372: data <= 8'h00;
	373: data <= 8'h30;
	374: data <= 8'h30;
	375: data <= 8'h00;
	// char 47, '/'
	376: data <= 8'h00;
	377: data <= 8'h04;
	378: data <= 8'h08;
	379: data <= 8'h10;
	380: data <= 8'h20;
	381: data <= 8'h40;
	382: data <= 8'h00;
	383: data <= 8'h00;
	// char 48, '0'
	384: data <= 8'h38;
	385: data <= 8'h44;
	386: data <= 8'h4c;
	387: data <= 8'h54;
	388: data <= 8'h64;
	389: data <= 8'h44;
	390: data <= 8'h38;
	391: data <= 8'h00;
	// char 49, '1'
	392: data <= 8'h10;
	393: data <= 8'h30;
	394: data <= 8'h10;
	395: data <= 8'h10;
	396: data <= 8'h10;
	397: data <= 8'h10;
	398: data <= 8'h38;
	399: data <= 8'h00;
	// char 50, '2'
	400: data <= 8'h38;
	401: data <= 8'h44;
	402: data <= 8'h04;
	403: data <= 8'h18;
	404: data <= 8'h20;
	405: data <= 8'h40;
	406: data <= 8'h7c;
	407: data <= 8'h00;
	// char 51, '3'
	408: data <= 8'h38;
	409: data <= 8'h44;
	410: data <= 8'h04;
	411: data <= 8'h38;
	412: data <= 8'h04;
	413: data <= 8'h44;
	414: data <= 8'h38;
	415: data <= 8'h00;
	// char 52, '4'
	416: data <= 8'h08;
	417: data <= 8'h18;
	418: data <= 8'h28;
	419: data <= 8'h48;
	420: data <= 8'h7c;
	421: data <= 8'h08;
	422: data <= 8'h08;
	423: data <= 8'h00;
	// char 53, '5'
	424: data <= 8'h7c;
	425: data <= 8'h40;
	426: data <= 8'h40;
	427: data <= 8'h78;
	428: data <= 8'h04;
	429: data <= 8'h44;
	430: data <= 8'h38;
	431: data <= 8'h00;
	// char 54, '6'
	432: data <= 8'h18;
	433: data <= 8'h20;
	434: data <= 8'h40;
	435: data <= 8'h78;
	436: data <= 8'h44;
	437: data <= 8'h44;
	438: data <= 8'h38;
	439: data <= 8'h00;
	// char 55, '7'
	440: data <= 8'h7c;
	441: data <= 8'h04;
	442: data <= 8'h08;
	443: data <= 8'h10;
	444: data <= 8'h20;
	445: data <= 8'h20;
	446: data <= 8'h20;
	447: data <= 8'h00;
	// char 56, '8'
	448: data <= 8'h38;
	449: data <= 8'h44;
	450: data <= 8'h44;
	451: data <= 8'h38;
	452: data <= 8'h44;
	453: data <= 8'h44;
	454: data <= 8'h38;
	455: data <= 8'h00;
	// char 57, '9'
	456: data <= 8'h38;
	457: data <= 8'h44;
	458: data <= 8'h44;
	459: data <= 8'h3c;
	460: data <= 8'h04;
	461: data <= 8'h08;
	462: data <= 8'h30;
	463: data <= 8'h00;
	// char 58, ':'
	464: data <= 8'h00;
	465: data <= 8'h00;
	466: data <= 8'h30;
	467: data <= 8'h30;
	468: data <= 8'h00;
	469: data <= 8'h30;
	470: data <= 8'h30;
	471: data <= 8'h00;
	// char 59, ';'
	472: data <= 8'h00;
	473: data <= 8'h00;
	474: data <= 8'h30;
	475: data <= 8'h30;
	476: data <= 8'h00;
	477: data <= 8'h30;
	478: data <= 8'h30;
	479: data <= 8'h20;
	// char 60, '<'
	480: data <= 8'h08;
	481: data <= 8'h10;
	482: data <= 8'h20;
	483: data <= 8'h40;
	484: data <= 8'h20;
	485: data <= 8'h10;
	486: data <= 8'h08;
	487: data <= 8'h00;
	// char 61, '='
	488: data <= 8'h00;
	489: data <= 8'h00;
	490: data <= 8'h7c;
	491: data <= 8'h00;
	492: data <= 8'h00;
	493: data <= 8'h7c;
	494: data <= 8'h00;
	495: data <= 8'h00;
	// char 62, '>'
	496: data <= 8'h20;
	497: data <= 8'h10;
	498: data <= 8'h08;
	499: data <= 8'h04;
	500: data <= 8'h08;
	501: data <= 8'h10;
	502: data <= 8'h20;
	503: data <= 8'h00;
	// char 63, '?'
	504: data <= 8'h38;
	505: data <= 8'h44;
	506: data <= 8'h04;
	507: data <= 8'h18;
	508: data <= 8'h10;
	509: data <= 8'h00;
	510: data <= 8'h10;
	511: data <= 8'h00;
	// char 64, '@'
	512: data <= 8'h38;
	513: data <= 8'h44;
	514: data <= 8'h5c;
	515: data <= 8'h54;
	516: data <= 8'h5c;
	517: data <= 8'h40;
	518: data <= 8'h38;
	519: data <= 8'h00;
	// char 65, 'A'
	520: data <= 8'h38;
	521: data <= 8'h44;
	522: data <= 8'h44;
	523: data <= 8'h44;
	524: data <= 8'h7c;
	525: data <= 8'h44;
	526: data <= 8'h44;
	527: data <= 8'h00;
	// char 66, 'B'
	528: data <= 8'h78;
	529: data <= 8'h44;
	530: data <= 8'h44;
	531: data <= 8'h78;
	532: data <= 8'h44;
	533: data <= 8'h44;
	534: data <= 8'h78;
	535: data <= 8'h00;
	// char 67, 'C'
	536: data <= 8'h38;
	537: data <= 8'h44;
	538: data <= 8'h40;
	539: data <= 8'h40;
	540: data <= 8'h40;
	541: data <= 8'h44;
	542: data <= 8'h38;
	543: data <= 8'h00;
	// char 68, 'D'
	544: data <= 8'h78;
	545: data <= 8'h44;
	546: data <= 8'h44;
	547: data <= 8'h44;
	548: data <= 8'h44;
	549: data <= 8'h44;
	550: data <= 8'h78;
	551: data <= 8'h00;
	// char 69, 'E'
	552: data <= 8'h7c;
	553: data <= 8'h40;
	554: data <= 8'h40;
	555: data <= 8'h78;
	556: data <= 8'h40;
	557: data <= 8'h40;
	558: data <= 8'h7c;
	559: data <= 8'h00;
	// char 70, 'F'
	560: data <= 8'h7c;
	561: data <= 8'h40;
	562: data <= 8'h40;
	563: data <= 8'h78;
	564: data <= 8'h40;
	565: data <= 8'h40;
	566: data <= 8'h40;
	567: data <= 8'h00;
	// char 71, 'G'
	568: data <= 8'h38;
	569: data <= 8'h44;
	570: data <= 8'h40;
	571: data <= 8'h5c;
	572: data <= 8'h44;
	573: data <= 8'h44;
	574: data <= 8'h3c;
	575: data <= 8'h00;
	// char 72, 'H'
	576: data <= 8'h44;
	577: data <= 8'h44;
	578: data <= 8'h44;
	579: data <= 8'h7c;
	580: data <= 8'h44;
	581: data <= 8'h44;
	582: data <= 8'h44;
	583: data <= 8'h00;
	// char 73, 'I'
	584: data <= 8'h38;
	585: data <= 8'h10;
	586: data <= 8'h10;
	587: data <= 8'h10;
	588: data <= 8'h10;
	589: data <= 8'h10;
	590: data <= 8'h38;
	591: data <= 8'h00;
	// char 74, 'J'
	592: data <= 8'h04;
	593: data <= 8'h04;
	594: data <= 8'h04;
	595: data <= 8'h04;
	596: data <= 8'h44;
	597: data <= 8'h44;
	598: data <= 8'h38;
	599: data <= 8'h00;
	// char 75, 'K'
	600: data <= 8'h44;
	601: data <= 8'h48;
	602: data <= 8'h50;
	603: data <= 8'h60;
	604: data <= 8'h50;
	605: data <= 8'h48;
	606: data <= 8'h44;
	607: data <= 8'h00;
	// char 76, 'L'
	608: data <= 8'h40;
	609: data <= 8'h40;
	610: data <= 8'h40;
	611: data <= 8'h40;
	612: data <= 8'h40;
	613: data <= 8'h40;
	614: data <= 8'h7c;
	615: data <= 8'h00;
	// char 77, 'M'
	616: data <= 8'h44;
	617: data <= 8'h6c;
	618: data <= 8'h54;
	619: data <= 8'h44;
	620: data <= 8'h44;
	621: data <= 8'h44;
	622: data <= 8'h44;
	623: data <= 8'h00;
	// char 78, 'N'
	624: data <= 8'h44;
	625: data <= 8'h64;
	626: data <= 8'h54;
	627: data <= 8'h4c;
	628: data <= 8'h44;
	629: data <= 8'h44;
	630: data <= 8'h44;
	631: data <= 8'h00;
	// char 79, 'O'
	632: data <= 8'h38;
	633: data <= 8'h44;
	634: data <= 8'h44;
	635: data <= 8'h44;
	636: data <= 8'h44;
	637: data <= 8'h44;
	638: data <= 8'h38;
	639: data <= 8'h00;
	// char 80, 'P'
	640: data <= 8'h78;
	641: data <= 8'h44;
	642: data <= 8'h44;
	643: data <= 8'h78;
	644: data <= 8'h40;
	645: data <= 8'h40;
	646: data <= 8'h40;
	647: data <= 8'h00;
	// char 81, 'Q'
	648: data <= 8'h38;
	649: data <= 8'h44;
	650: data <= 8'h44;
	651: data <= 8'h44;
	652: data <= 8'h54;
	653: data <= 8'h48;
	654: data <= 8'h34;
	655: data <= 8'h00;
	// char 82, 'R'
	656: data <= 8'h78;
	657: data <= 8'h44;
	658: data <= 8'h44;
	659: data <= 8'h78;
	660: data <= 8'h48;
	661: data <= 8'h44;
	662: data <= 8'h44;
	663: data <= 8'h00;
	// char 83, 'S'
	664: data <= 8'h38;
	665: data <= 8'h44;
	666: data <= 8'h40;
	667: data <= 8'h38;
	668: data <= 8'h04;
	669: data <= 8'h44;
	670: data <= 8'h38;
	671: data <= 8'h00;
	// char 84, 'T'
	672: data <= 8'h7c;
	673: data <= 8'h10;
	674: data <= 8'h10;
	675: data <= 8'h10;
	676: data <= 8'h10;
	677: data <= 8'h10;
	678: data <= 8'h10;
	679: data <= 8'h00;
	// char 85, 'U'
	680: data <= 8'h44;
	681: data <= 8'h44;
	682: data <= 8'h44;
	683: data <= 8'h44;
	684: data <= 8'h44;
	685: data <= 8'h44;
	686: data <= 8'h38;
	687: data <= 8'h00;
	// char 86, 'V'
	688: data <= 8'h44;
	689: data <= 8'h44;
	690: data <= 8'h44;
	691: data <= 8'h44;
	692: data <= 8'h44;
	693: data <= 8'h28;
	694: data <= 8'h10;
	695: data <= 8'h00;
	// char 87, 'W'
	696: data <= 8'h44;
	697: data <= 8'h44;
	698: data <= 8'h54;
	699: data <= 8'h54;
	700: data <= 8'h54;
	701: data <= 8'h54;
	702: data <= 8'h28;
	703: data <= 8'h00;
	// char 88, 'X'
	704: data <= 8'h44;
	705: data <= 8'h44;
	706: data <= 8'h28;
	707: data <= 8'h10;
	708: data <= 8'h28;
	709: data <= 8'h44;
	710: data <= 8'h44;
	711: data <= 8'h00;
	// char 89, 'Y'
	712: data <= 8'h44;
	713: data <= 8'h44;
	714: data <= 8'h44;
	715: data <= 8'h28;
	716: data <= 8'h10;
	717: data <= 8'h10;
	718: data <= 8'h10;
	719: data <= 8'h00;
	// char 90, 'Z'
	720: data <= 8'h78;
	721: data <= 8'h08;
	722: data <= 8'h10;
	723: data <= 8'h20;
	724: data <= 8'h40;
	725: data <= 8'h40;
	726: data <= 8'h78;
	727: data <= 8'h00;
	// char 91, '['
	728: data <= 8'h38;
	729: data <= 8'h20;
	730: data <= 8'h20;
	731: data <= 8'h20;
	732: data <= 8'h20;
	733: data <= 8'h20;
	734: data <= 8'h38;
	735: data <= 8'h00;
	// char 92, '\'
	736: data <= 8'h00;
	737: data <= 8'h40;
	738: data <= 8'h20;
	739: data <= 8'h10;
	740: data <= 8'h08;
	741: data <= 8'h04;
	742: data <= 8'h00;
	743: data <= 8'h00;
	// char 93, ']'
	744: data <= 8'h38;
	745: data <= 8'h08;
	746: data <= 8'h08;
	747: data <= 8'h08;
	748: data <= 8'h08;
	749: data <= 8'h08;
	750: data <= 8'h38;
	751: data <= 8'h00;
	// char 94, '^'
	752: data <= 8'h10;
	753: data <= 8'h28;
	754: data <= 8'h44;
	755: data <= 8'h00;
	756: data <= 8'h00;
	757: data <= 8'h00;
	758: data <= 8'h00;
	759: data <= 8'h00;
	// char 95, '_'
	760: data <= 8'h00;
	761: data <= 8'h00;
	762: data <= 8'h00;
	763: data <= 8'h00;
	764: data <= 8'h00;
	765: data <= 8'h00;
	766: data <= 8'h00;
	767: data <= 8'hfc;
	// char 96, '`'
	768: data <= 8'h30;
	769: data <= 8'h30;
	770: data <= 8'h10;
	771: data <= 8'h00;
	772: data <= 8'h00;
	773: data <= 8'h00;
	774: data <= 8'h00;
	775: data <= 8'h00;
	// char 97, 'a'
	776: data <= 8'h00;
	777: data <= 8'h00;
	778: data <= 8'h38;
	779: data <= 8'h04;
	780: data <= 8'h3c;
	781: data <= 8'h44;
	782: data <= 8'h3c;
	783: data <= 8'h00;
	// char 98, 'b'
	784: data <= 8'h40;
	785: data <= 8'h40;
	786: data <= 8'h78;
	787: data <= 8'h44;
	788: data <= 8'h44;
	789: data <= 8'h44;
	790: data <= 8'h78;
	791: data <= 8'h00;
	// char 99, 'c'
	792: data <= 8'h00;
	793: data <= 8'h00;
	794: data <= 8'h38;
	795: data <= 8'h44;
	796: data <= 8'h40;
	797: data <= 8'h44;
	798: data <= 8'h38;
	799: data <= 8'h00;
	// char 100, 'd'
	800: data <= 8'h04;
	801: data <= 8'h04;
	802: data <= 8'h3c;
	803: data <= 8'h44;
	804: data <= 8'h44;
	805: data <= 8'h44;
	806: data <= 8'h3c;
	807: data <= 8'h00;
	// char 101, 'e'
	808: data <= 8'h00;
	809: data <= 8'h00;
	810: data <= 8'h38;
	811: data <= 8'h44;
	812: data <= 8'h78;
	813: data <= 8'h40;
	814: data <= 8'h38;
	815: data <= 8'h00;
	// char 102, 'f'
	816: data <= 8'h18;
	817: data <= 8'h20;
	818: data <= 8'h20;
	819: data <= 8'h78;
	820: data <= 8'h20;
	821: data <= 8'h20;
	822: data <= 8'h20;
	823: data <= 8'h00;
	// char 103, 'g'
	824: data <= 8'h00;
	825: data <= 8'h00;
	826: data <= 8'h3c;
	827: data <= 8'h44;
	828: data <= 8'h44;
	829: data <= 8'h3c;
	830: data <= 8'h04;
	831: data <= 8'h38;
	// char 104, 'h'
	832: data <= 8'h40;
	833: data <= 8'h40;
	834: data <= 8'h70;
	835: data <= 8'h48;
	836: data <= 8'h48;
	837: data <= 8'h48;
	838: data <= 8'h48;
	839: data <= 8'h00;
	// char 105, 'i'
	840: data <= 8'h10;
	841: data <= 8'h00;
	842: data <= 8'h10;
	843: data <= 8'h10;
	844: data <= 8'h10;
	845: data <= 8'h10;
	846: data <= 8'h18;
	847: data <= 8'h00;
	// char 106, 'j'
	848: data <= 8'h08;
	849: data <= 8'h00;
	850: data <= 8'h18;
	851: data <= 8'h08;
	852: data <= 8'h08;
	853: data <= 8'h08;
	854: data <= 8'h48;
	855: data <= 8'h30;
	// char 107, 'k'
	856: data <= 8'h40;
	857: data <= 8'h40;
	858: data <= 8'h48;
	859: data <= 8'h50;
	860: data <= 8'h60;
	861: data <= 8'h50;
	862: data <= 8'h48;
	863: data <= 8'h00;
	// char 108, 'l'
	864: data <= 8'h10;
	865: data <= 8'h10;
	866: data <= 8'h10;
	867: data <= 8'h10;
	868: data <= 8'h10;
	869: data <= 8'h10;
	870: data <= 8'h18;
	871: data <= 8'h00;
	// char 109, 'm'
	872: data <= 8'h00;
	873: data <= 8'h00;
	874: data <= 8'h68;
	875: data <= 8'h54;
	876: data <= 8'h54;
	877: data <= 8'h44;
	878: data <= 8'h44;
	879: data <= 8'h00;
	// char 110, 'n'
	880: data <= 8'h00;
	881: data <= 8'h00;
	882: data <= 8'h70;
	883: data <= 8'h48;
	884: data <= 8'h48;
	885: data <= 8'h48;
	886: data <= 8'h48;
	887: data <= 8'h00;
	// char 111, 'o'
	888: data <= 8'h00;
	889: data <= 8'h00;
	890: data <= 8'h38;
	891: data <= 8'h44;
	892: data <= 8'h44;
	893: data <= 8'h44;
	894: data <= 8'h38;
	895: data <= 8'h00;
	// char 112, 'p'
	896: data <= 8'h00;
	897: data <= 8'h00;
	898: data <= 8'h78;
	899: data <= 8'h44;
	900: data <= 8'h44;
	901: data <= 8'h44;
	902: data <= 8'h78;
	903: data <= 8'h40;
	// char 113, 'q'
	904: data <= 8'h00;
	905: data <= 8'h00;
	906: data <= 8'h3c;
	907: data <= 8'h44;
	908: data <= 8'h44;
	909: data <= 8'h44;
	910: data <= 8'h3c;
	911: data <= 8'h04;
	// char 114, 'r'
	912: data <= 8'h00;
	913: data <= 8'h00;
	914: data <= 8'h58;
	915: data <= 8'h24;
	916: data <= 8'h20;
	917: data <= 8'h20;
	918: data <= 8'h70;
	919: data <= 8'h00;
	// char 115, 's'
	920: data <= 8'h00;
	921: data <= 8'h00;
	922: data <= 8'h38;
	923: data <= 8'h40;
	924: data <= 8'h38;
	925: data <= 8'h04;
	926: data <= 8'h38;
	927: data <= 8'h00;
	// char 116, 't'
	928: data <= 8'h00;
	929: data <= 8'h20;
	930: data <= 8'h78;
	931: data <= 8'h20;
	932: data <= 8'h20;
	933: data <= 8'h28;
	934: data <= 8'h10;
	935: data <= 8'h00;
	// char 117, 'u'
	936: data <= 8'h00;
	937: data <= 8'h00;
	938: data <= 8'h48;
	939: data <= 8'h48;
	940: data <= 8'h48;
	941: data <= 8'h58;
	942: data <= 8'h28;
	943: data <= 8'h00;
	// char 118, 'v'
	944: data <= 8'h00;
	945: data <= 8'h00;
	946: data <= 8'h44;
	947: data <= 8'h44;
	948: data <= 8'h44;
	949: data <= 8'h28;
	950: data <= 8'h10;
	951: data <= 8'h00;
	// char 119, 'w'
	952: data <= 8'h00;
	953: data <= 8'h00;
	954: data <= 8'h44;
	955: data <= 8'h44;
	956: data <= 8'h54;
	957: data <= 8'h7c;
	958: data <= 8'h28;
	959: data <= 8'h00;
	// char 120, 'x'
	960: data <= 8'h00;
	961: data <= 8'h00;
	962: data <= 8'h48;
	963: data <= 8'h48;
	964: data <= 8'h30;
	965: data <= 8'h48;
	966: data <= 8'h48;
	967: data <= 8'h00;
	// char 121, 'y'
	968: data <= 8'h00;
	969: data <= 8'h00;
	970: data <= 8'h48;
	971: data <= 8'h48;
	972: data <= 8'h48;
	973: data <= 8'h38;
	974: data <= 8'h10;
	975: data <= 8'h60;
	// char 122, 'z'
	976: data <= 8'h00;
	977: data <= 8'h00;
	978: data <= 8'h78;
	979: data <= 8'h08;
	980: data <= 8'h30;
	981: data <= 8'h40;
	982: data <= 8'h78;
	983: data <= 8'h00;
	// char 123, '{'
	984: data <= 8'h18;
	985: data <= 8'h20;
	986: data <= 8'h20;
	987: data <= 8'h60;
	988: data <= 8'h20;
	989: data <= 8'h20;
	990: data <= 8'h18;
	991: data <= 8'h00;
	// char 124, '|'
	992: data <= 8'h10;
	993: data <= 8'h10;
	994: data <= 8'h10;
	995: data <= 8'h00;
	996: data <= 8'h10;
	997: data <= 8'h10;
	998: data <= 8'h10;
	999: data <= 8'h00;
	// char 125, '}'
	1000: data <= 8'h30;
	1001: data <= 8'h08;
	1002: data <= 8'h08;
	1003: data <= 8'h0c;
	1004: data <= 8'h08;
	1005: data <= 8'h08;
	1006: data <= 8'h30;
	1007: data <= 8'h00;
	// char 126, '~'
	1008: data <= 8'h28;
	1009: data <= 8'h50;
	1010: data <= 8'h00;
	1011: data <= 8'h00;
	1012: data <= 8'h00;
	1013: data <= 8'h00;
	1014: data <= 8'h00;
	1015: data <= 8'h00;
	// char 127, '.'
	1016: data <= 8'h00;
	1017: data <= 8'h00;
	1018: data <= 8'h00;
	1019: data <= 8'h00;
	1020: data <= 8'h00;
	1021: data <= 8'h00;
	1022: data <= 8'h00;
	1023: data <= 8'h00;

//       10'h000: data <= 8'h00;
       default: data <= 8'h00;
     endcase

endmodule
