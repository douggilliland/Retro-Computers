-- PDP-11/70 build
--
--	http://land-boards.com/blwiki/index.php?title=PDP-11_ON_RETRO-EP4CE15
-- Wiki page: http://land-boards.com/blwiki/index.php?title=PDP-11_ON_RETRO-EP4CE15
--	Front Panel: 
--	Hackaday page - https://hackaday.io/project/179642-pdp-11-on-a-fpga
--
-- Copyright (c) 2008-2021 Sytse van Slooten
--
-- Permission is hereby granted to any person obtaining a copy of these VHDL source files and
-- other language source files and associated documentation files ("the materials") to use
-- these materials solely for personal, non-commercial purposes.
-- You are also granted permission to make changes to the materials, on the condition that this
-- copyright notice is retained unchanged.
--
-- The materials are distributed in the hope that they will be useful, but WITHOUT ANY WARRANTY;
-- without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
--

-- $Revision$

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
--use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;

entity top is
   port(
      clkin 		: in std_logic;

		-- Switches and PEDs
		i_SS			: in std_logic_vector(8 downto 1);
		i_PB			: in std_logic_vector(8 downto 1);
		o_LED			: OUT std_logic_vector(8 downto 1);
		
		-- VGA (2:2:2)
      vgar			: out std_logic_vector(1 downto 0);
      vgag			: out std_logic_vector(1 downto 0);
      vgab			: out std_logic_vector(1 downto 0);
      vgah			: out std_logic;
      vgav			: out std_logic;

		-- PS/2 keyboard
      ps2k_c		: in std_logic;
      ps2k_d		: in std_logic;

		-- Serial port
		-- USB-to-Serial - 9600/8/n/1 debug output from microcode
      tx1			: out std_logic;
      rx1			: in std_logic;
      rts1			: out std_logic;
      cts1			: in std_logic;

		-- SD card
      sdcard_cs	: out std_logic;
      sdcard_mosi : out std_logic;
      sdcard_sclk : out std_logic;
      sdcard_miso : in std_logic;

		-- Ethernet, enc424j600 controller interface
      xu_cs			: out std_logic;
      xu_mosi		: out std_logic;
      xu_sclk		: out std_logic;
      xu_miso		: in std_logic;
      xu_debug_tx	: out std_logic;

		-- Uses the SDRAM as the main storage space
      dram_addr	: out std_logic_vector(12 downto 0);
      dram_dq		: inout std_logic_vector(15 downto 0);
      dram_ba_1	: out std_logic;
      dram_ba_0	: out std_logic;
      dram_udqm	: out std_logic;
      dram_ldqm	: out std_logic;
      dram_ras_n	: out std_logic;
      dram_cas_n	: out std_logic;
      dram_cke		: out std_logic;
      dram_clk		: out std_logic;
      dram_we_n	: out std_logic;
      dram_cs_n	: out std_logic
   );
end top;

architecture implementation of top is

component unibus is
   port(
-- clocks and reset
      clk : in std_logic;													-- cpu clock
      clk50mhz : in std_logic;											-- 50Mhz clock for peripherals
      reset : in std_logic;												-- active '1' synchronous reset
		
-- bus interface
      addr				: out std_logic_vector(21 downto 0);		-- physical address driven out to the bus by cpu or busmaster peripherals
      dati				: in std_logic_vector(15 downto 0);			-- data input to cpu or busmaster peripherals
      dato				: out std_logic_vector(15 downto 0);		-- data output from cpu or busmaster peripherals
      control_dati	: out std_logic;									-- if '1', this is an input cycle
      control_dato	: out std_logic;									-- if '1', this is an output cycle
      control_datob	: out std_logic;									-- if '1', the current output cycle is for a byte
      addr_match		: in std_logic;									-- '1' if the address is recognized

-- debug & blinkenlights
      ifetch			: out std_logic;									-- '1' if this cycle is an ifetch cycle
      iwait				: out std_logic;									-- '1' if the cpu is in wait state
      cpu_addr_v		: out std_logic_vector(15 downto 0);		-- virtual address from cpu, for debug and general interest

-- rl controller
      have_rl				: in integer range 0 to 1 := 0;			-- enable conditional compilation
      rl_sdcard_cs		: out std_logic;
      rl_sdcard_mosi		: out std_logic;
      rl_sdcard_sclk		: out std_logic;
      rl_sdcard_miso		: in std_logic := '0';
      rl_sdcard_debug	: out std_logic_vector(3 downto 0);		-- debug/blinkenlights

-- rk controller
      have_rk				: in integer range 0 to 1 := 0;				-- enable conditional compilation
      have_rk_num			: in integer range 1 to 8 := 8;				-- active number of drives on the controller; set to < 8 to save core
      rk_sdcard_cs		: out std_logic;
      rk_sdcard_mosi 	: out std_logic;
      rk_sdcard_sclk 	: out std_logic;
      rk_sdcard_miso 	: in std_logic := '0';
      rk_sdcard_debug	: out std_logic_vector(3 downto 0);		-- debug/blinkenlights

-- rh controller
      have_rh				: in integer range 0 to 1 := 0;				-- enable conditional compilation
      rh_sdcard_cs		: out std_logic;
      rh_sdcard_mosi 	: out std_logic;
      rh_sdcard_sclk 	: out std_logic;
      rh_sdcard_miso 	: in std_logic := '0';
      rh_sdcard_debug	: out std_logic_vector(3 downto 0);		-- debug/blinkenlights
      rh_type				: in integer range 4 to 7 := 6;

-- xu enc424j600 controller interface
      have_xu			: in integer range 0 to 1 := 0;				-- enable conditional compilation
      have_xu_debug	: in integer range 0 to 1 := 1;				-- enable debug core
      xu_cs				: out std_logic;
      xu_mosi			: out std_logic;
      xu_sclk			: out std_logic;
      xu_miso			: in std_logic := '0';
      xu_debug_tx		: out std_logic;

-- kl11, console ports
-- rs232, 9600/8/n/1 debug output from microcode
      have_kl11		: in integer range 0 to 4 := 4;				-- conditional compilation - number of kl11 controllers to include. Should normally be at least 1

      tx0				: out std_logic;
      rx0				: in std_logic := '1';
      rts0				: out std_logic;
      cts0				: in std_logic := '0';
      kl0_bps			: in integer range 1200 to 230400 := 9600;	-- bps rate - don't set over 38400 for interrupt control applications
      kl0_force7bit	: in integer range 0 to 1 := 1;					-- zero out high order bit on transmission and reception
      kl0_rtscts		: in integer range 0 to 1 := 1;					-- conditional compilation switch for rts and cts signals; also implies to include core that implements a silo buffer

      tx1				: out std_logic;
      rx1 				: in std_logic := '1';
      rts1				: out std_logic;
      cts1				: in std_logic := '0';
      kl1_bps			: in integer range 1200 to 230400 := 9600;
      kl1_force7bit	: in integer range 0 to 1 := 1;
      kl1_rtscts		: in integer range 0 to 1 := 0;

      tx2				: out std_logic;
      rx2				: in std_logic := '1';
      rts2				: out std_logic;
      cts2				: in std_logic := '0';
      kl2_bps			: in integer range 1200 to 230400 := 9600;
      kl2_force7bit	: in integer range 0 to 1 := 1;
      kl2_rtscts		: in integer range 0 to 1 := 0;

      tx3				: out std_logic;
      rx3				: in std_logic := '1';
      rts3				: out std_logic;
      cts3				: in std_logic := '0';
      kl3_bps			: in integer range 1200 to 230400 := 9600;
      kl3_force7bit	: in integer range 0 to 1 := 1;
      kl3_rtscts		: in integer range 0 to 1 := 0;

-- dr11c, universal interface

      have_dr11c						: in integer range 0 to 1 := 0;		-- conditional compilation
      have_dr11c_loopback			: in integer range 0 to 1 := 0;		-- for testing only - zdrc
      have_dr11c_signal_stretch	: in integer range 0 to 127 := 7;	-- the signals ndr*, dxm, init will be stretched to this many cpu cycles

      dr11c_in		: in std_logic_vector(15 downto 0) := (others => '0');
      dr11c_out	: out std_logic_vector(15 downto 0);
      dr11c_reqa	: in std_logic := '0';
      dr11c_reqb	: in std_logic := '0';
      dr11c_csr0	: out std_logic;
      dr11c_csr1	: out std_logic;
      dr11c_ndr	: out std_logic;                                     -- new data ready : dr11c_out has new data
      dr11c_ndrlo	: out std_logic;                                   -- new data ready : dr11c_out(7 downto 0) has new data
      dr11c_ndrhi	: out std_logic;                                   -- new data ready : dr11c_out(15 downto 8) has new data
      dr11c_dxm	: out std_logic;                                     -- data transmitted : dr11c_in data has been read by the cpu
      dr11c_init	: out std_logic;                                    -- unibus reset propagated out to the user device

-- minc-11

      have_mncad			: in integer range 0 to 1 := 0;                     	-- mncad: a/d, max one card in a system
      have_mnckw			: in integer range 0 to 2 := 0;                     	-- mnckw: clock, either one or two
      have_mncaa			: in integer range 0 to 1 := 0;                     	-- mncaa: d/a
      have_mncdi			: in integer range 0 to 1 := 0;                     	-- mncdo: digital in
      have_mncdo			: in integer range 0 to 1 := 0;                     	-- mncdo: digital out
      ad_start				: out std_logic;                                      -- interface from mncad to a/d hardware : '1' signals to start converting
      ad_done				: in std_logic := '1';                                -- interface from mncad to a/d hardware : '1' signals to the mncad that the a/d has completed a conversion
      ad_channel			: out std_logic_vector(5 downto 0);                 	-- interface from mncad to a/d hardware : the channel number for the current command
      ad_nxc				: in std_logic := '1';                                -- interface from mncad to a/d hardware : '1' signals to the mncad that the required channel does not exist
      ad_sample			: in std_logic_vector(11 downto 0) := "000000000000";	-- interface from mncad to a/d hardware : the value of the last sample
      kw_st1in				: in std_logic := '0';                                -- mnckw0 st1 signal input, active on rising edge
      kw_st2in				: in std_logic := '0';                                -- mnckw0 st2 signal input, active on rising edge
      kw_st1out			: out std_logic;                                     	-- mnckw0 st1 output pulse (actually : copy of the st1flag in the csr
      kw_st2out			: out std_logic;                                     	-- mnckw0 st2 output pulse
      kw_clkov				: out std_logic;                                      -- mnckw0 clkovf output pulse
      da_dac1				: out std_logic_vector(11 downto 0);
      da_dac2				: out std_logic_vector(11 downto 0);
      da_dac3				: out std_logic_vector(11 downto 0);
      da_dac4				: out std_logic_vector(11 downto 0);
      have_diloopback	: in integer range 0 to 1 := 0;                					-- set to 1 to loop back mncdo0 to mncdi0 internally for testing
      di_dir				: in std_logic_vector(15 downto 0) := "0000000000000000";   -- mncdi0 data input register
      di_strobe			: in std_logic := '0';
      di_reply				: out std_logic;
      di_pgmout			: out std_logic;
      di_event				: out std_logic;
      do_dor				: out std_logic_vector(15 downto 0);
      do_hb_strobe		: out std_logic;
      do_lb_strobe		: out std_logic;
      do_reply				: in std_logic := '0';

-- cpu console, switches and display register
      have_csdr : in integer range 0 to 1 := 1;

-- clock
      have_kw11l : in integer range 0 to 1 := 1;			-- conditional compilation
      kw11l_hz : in integer range 50 to 800 := 60;			-- valid values are 50, 60, 800

-- model code
      modelcode	: in integer range 0 to 255;				-- mostly used are 20,34,44,45,70,94; others are less well tested
      have_fp		: in integer range 0 to 2 := 2;			-- fp11 switch; 0=don't include; 1=include; 2=include if the cpu model can support fp11
      have_fpa		: in integer range 0 to 1 := 1;			-- floating point accelerator present with J11 cpu

-- cpu initial r7 and psw
      init_r7 : in std_logic_vector(15 downto 0) := x"ea10";	-- start address after reset f600 = o'173000' = m9312 hi rom; ea10 = 165020 = m9312 lo rom
      init_psw : in std_logic_vector(15 downto 0) := x"00e0";	-- initial psw for kernel mode, primary register set, priority 7

-- console
      cons_load		: in std_logic := '0';
      cons_exa			: in std_logic := '0';									-- Examine memory
      cons_dep			: in std_logic := '0';									-- Deposit
      cons_cont		: in std_logic := '0';									-- continue, pulse '1'
      cons_ena			: in std_logic := '1';									-- ena/halt, '1' is enable
      cons_start		: in std_logic := '0';
      cons_sw			: in std_logic_vector(21 downto 0) := (others => '0');
      cons_adss_mode : in std_logic_vector(1 downto 0) := (others => '0');
      cons_adss_id	: in std_logic := '0';
      cons_adss_cons : in std_logic := '0';
      cons_consphy	: out std_logic_vector(21 downto 0);
      cons_progphy	: out std_logic_vector(21 downto 0);
      cons_br			: out std_logic_vector(15 downto 0);
      cons_shfr		: out std_logic_vector(15 downto 0);
      cons_maddr		: out std_logic_vector(15 downto 0);				-- microcode address fpu/cpu
      cons_dr			: out std_logic_vector(15 downto 0);
      cons_parh		: out std_logic;
      cons_parl		: out std_logic;

      cons_adrserr	: out std_logic;
      cons_run			: out std_logic;		-- '1' if executing instructions (incl wait)
      cons_pause		: out std_logic;		-- '1' if bus has been relinquished to npr
      cons_master		: out std_logic;		-- '1' if cpu is bus master and not running
      cons_kernel		: out std_logic;		-- '1' if kernel mode
      cons_super		: out std_logic;		-- '1' if super mode
      cons_user		: out std_logic;		-- '1' if user mode
      cons_id			: out std_logic;		-- '0' if instruction, '1' if data AND data mapping is enabled in the mmu
      cons_map16		: out std_logic;		-- '1' if 16-bit mapping
      cons_map18		: out std_logic;		-- '1' if 18-bit mapping
      cons_map22		: out std_logic		-- '1' if 22-bit mapping
   );
end component;

component vt is
   port(
      vga_hsync	: out std_logic;			-- horizontal sync
      vga_vsync	: out std_logic;			-- vertical sync
      vga_fb		: out std_logic;			-- output - full
      vga_ht		: out std_logic;			-- output - half

-- serial port
      tx				: out std_logic;										-- transmit
      rx				: in std_logic;										-- receive
      rts			: out std_logic;										-- request to send
      cts			: in std_logic := '0';								-- clear to send
      bps			: in integer range 1200 to 230400 := 9600;	-- bps rate - don't set to more than 38400
      force7bit	: in integer range 0 to 1 := 0;					-- zero out high order bit on transmission and reception
      rtscts		: in integer range 0 to 1 := 0;					-- conditional compilation switch for rts and cts signals; also implies to include core that implements a silo buffer

-- ps2 keyboard
      ps2k_c : in std_logic;			-- clock
      ps2k_d : in std_logic;			-- data

-- debug & blinkenlights
      ifetch		: out std_logic;								-- ifetch : the cpu is running an instruction fetch cycle
      iwait			: out std_logic;								-- iwait : the cpu is in wait state
      teste			: in std_logic := '0';						-- teste : display 24*80 capital E without changing the display buffer
      testf			: in std_logic := '0';						-- testf : display 24*80 all pixels on
      vga_debug	: out std_logic_vector(15 downto 0);	-- debug output from microcode
      vga_bl		: out std_logic_vector(9 downto 0);		-- blinkenlight vector

-- vt type code : 100 or 105
      vttype				: in integer range 100 to 105 := 100;	-- vt100 or vt105
      vga_cursor_block	: in std_logic := '1';						-- cursor is block ('1') or underline ('0')
      vga_cursor_blink	: in std_logic := '1';						-- cursor blinks ('1') or not ('0')
      have_act_seconds	: in integer range 0 to 7200 := 1800;	-- auto screen off time, in seconds; 0 means disabled
      have_act				: in integer range 1 to 2 := 2;			-- auto screen off counter reset by keyboard and serial port activity (1) or keyboard only (2)

-- clock & reset
      cpuclk	: in std_logic;		-- cpuclk : should be around 10MHz, give or take a few
      clk50mhz	: in std_logic;		-- clk50mhz : used for vga signal timing
      reset		: in std_logic			-- reset
   );
end component;

component pll is
   port(
      inclk0	: in std_logic := '0';
      c0			: out std_logic
   );
end component;

signal c0 					: std_logic;

signal cpuclk 				: std_logic := '0';
signal cpureset			: std_logic := '1';
signal cpuresetlength	: integer range 0 to 63 := 63;
signal slowreset			: std_logic;
signal slowresetdelay	: integer range 0 to 4095 := 4095;
signal vtreset				: std_logic := '1';

signal ifetch				: std_logic;
signal iwait				: std_logic;
signal reset				: std_logic;
signal txtx0				: std_logic;
signal rxrx0				: std_logic;
signal txtx1				: std_logic;
signal rxrx1				: std_logic;
signal rtsrts1				: std_logic;
signal ctscts1				: std_logic;

signal addr				: std_logic_vector(21 downto 0);
signal addrq			: std_logic_vector(21 downto 0);
signal dati				: std_logic_vector(15 downto 0);
signal dato				: std_logic_vector(15 downto 0);
signal control_dati	: std_logic;
signal control_dato	: std_logic;
signal control_datob : std_logic;

signal have_rl			: integer range 0 to 1;
signal rl_cs			: std_logic;
signal rl_mosi			: std_logic;
signal rl_miso			: std_logic;
signal rl_sclk			: std_logic;
signal rl_sddebug		: std_logic_vector(3 downto 0);

signal have_rk			: integer range 0 to 1;
signal rk_cs			: std_logic;
signal rk_mosi			: std_logic;
signal rk_miso			: std_logic;
signal rk_sclk			: std_logic;
signal rk_sddebug		: std_logic_vector(3 downto 0);

signal have_rh			: integer range 0 to 1;
signal rh_cs			: std_logic;
signal rh_mosi			: std_logic;
signal rh_miso			: std_logic;
signal rh_sclk			: std_logic;
signal rh_sddebug		: std_logic_vector(3 downto 0);

signal have_kl11		: integer range 0 to 1;
signal have_xu			: integer range 0 to 1;

signal sddebug			: std_logic_vector(3 downto 0);

signal vga_hsync		: std_logic;
signal vga_vsync		: std_logic;
signal vga_fb			: std_logic;
signal vga_ht			: std_logic;

signal dram_match		: std_logic;
signal dram_counter	: integer range 0 to 32767;
signal dram_wait		: integer range 0 to 15;

signal resetbtn		: std_logic;
signal sw				: std_logic_vector(5 downto 0);
signal greenled		: std_logic_vector(4 downto 0);

type dram_fsm_type is (
   dram_init,
   dram_poweron,
   dram_pwron_pre, dram_pwron_prew,
   dram_pwron_ref, dram_pwron_refw,
   dram_pwron_mrs, dram_pwron_mrsw,
   dram_c1,
   dram_c2,
   dram_c3,
   dram_c4,
   dram_c5,
   dram_c6,
   dram_c7,
   dram_c8,
   dram_c9,
   dram_c10,
   dram_c11,
   dram_c12,
   dram_c13,
   dram_c14,
   dram_c15,
   dram_c16,
   dram_idle
);
signal dram_fsm : dram_fsm_type := dram_init;

begin

-- Mapping to SWITCHES-LEDS-2 Card

-- Pushbuttons (left to right)
resetbtn	<= i_PB(8);				-- CPU Reset button

-- Slide Switches (left to right)
sw(5)		<= i_SS(6);				-- Unused
sw(4)		<= i_SS(5);				-- unused
sw(3)		<= i_SS(4);				-- 1 = K11 Serial TTY present
sw(2)		<= not i_SS(3);		-- RH (RP) drive when on
sw(1)		<= not i_SS(2);		-- RK drive when on
sw(0)		<= not i_SS(1);		-- PL drive when on

-- LEDs (left to right)
o_LED(8) <= '1';					-- POWER LED
o_LED(7)	<= not greenled(1);	-- Off = SD card. On = SDHC card
o_LED(6) <= greenled(4);		-- Instruction Fetch
o_LED(5) <= greenled(3);		-- Write to SD Card?
o_LED(4)	<= greenled(2);		-- Read from SD card?
o_LED(3)	<= i_SS(3);				-- RH (RP) drive when on
o_LED(2)	<= i_SS(2);				-- RK drive when on
o_LED(1)	<= i_SS(1);				-- RL drive when on


   pll0: pll port map(
      inclk0 => clkin,
      c0 => c0
   );

--   c0 <= clkin;

   pdp11: unibus port map(

      modelcode => 70,

      reset				=> cpureset,
      clk50mhz			=> clkin,
      clk				=> cpuclk,
		
      addr				=> addr,
      dati				=> dati,
      dato				=> dato,
      control_dati	=> control_dati,
      control_dato	=> control_dato,
      control_datob	=> control_datob,
      addr_match		=> dram_match,

      ifetch			=> ifetch,
      iwait				=> iwait,

      have_rl				=> have_rl,
      rl_sdcard_cs		=> rl_cs,
      rl_sdcard_mosi 	=> rl_mosi,
      rl_sdcard_sclk 	=> rl_sclk,
      rl_sdcard_miso 	=> rl_miso,
      rl_sdcard_debug 	=> rl_sddebug,

      have_rk				=> have_rk,
      rk_sdcard_cs		=> rk_cs,
      rk_sdcard_mosi		=> rk_mosi,
      rk_sdcard_sclk		=> rk_sclk,
      rk_sdcard_miso		=> rk_miso,
      rk_sdcard_debug	=> rk_sddebug,

      have_rh				=> have_rh,
      rh_sdcard_cs		=> rh_cs,
      rh_sdcard_mosi		=> rh_mosi,
      rh_sdcard_sclk		=> rh_sclk,
      rh_sdcard_miso		=> rh_miso,
      rh_sdcard_debug	=> rh_sddebug,

      have_kl11			=> have_kl11,
      rx0					=> rxrx0,
      tx0					=> txtx0,
      rx1					=> rxrx1,
      tx1					=> txtx1,
		rts1					=> rtsrts1,
		cts1					=> ctscts1,

      have_xu				=> 0,			-- Not enough resources in a 5CEFA2 FPGA
      xu_cs					=> xu_cs,
      xu_mosi				=> xu_mosi,
      xu_sclk				=> xu_sclk,
      xu_miso				=> xu_miso,
      xu_debug_tx			=> xu_debug_tx
   );

   vt0: vt port map(
      vga_hsync			=> vga_hsync,
      vga_vsync			=> vga_vsync,
      vga_fb				=> vga_fb,
      vga_ht				=> vga_ht,

      rx						=> txtx0,
      tx						=> rxrx0,

      ps2k_c				=> ps2k_c,
      ps2k_d				=> ps2k_d,

      vttype => 100,

      cpuclk				=> cpuclk,
      clk50mhz				=> clkin,
      reset					=> vtreset
   );


   reset <= (not resetbtn) ; -- or power_on_reset;

   -- Status LEDs
	greenled<= ifetch & sddebug;

   -- Map to FPGA pins
	tx1 <= txtx1;
   rxrx1 <= rx1;
	rts1 <= rtsrts1;
	ctscts1 <= cts1;

   sddebug		<= rh_sddebug when have_rh = 1 else
						rl_sddebug when have_rl = 1 else
						rk_sddebug;
   sdcard_cs	<= rh_cs when have_rh = 1 else 
						rl_cs when have_rl = 1 else
						rk_cs;
   sdcard_mosi	<= rh_mosi when have_rh = 1 else 
						rl_mosi when have_rl = 1 else 
						rk_mosi;
   sdcard_sclk <= rh_sclk when have_rh = 1 else
						rl_sclk when have_rl = 1 else
						rk_sclk;
   rh_miso		<= sdcard_miso;
   rl_miso		<= sdcard_miso;
   rk_miso		<= sdcard_miso;

	-- The hexadecimal RGB code of Amber color is #FFBF00
   vgar <=	"11" when vga_fb = '1' else
				"10" when vga_ht = '1' else
				"00";
   vgag <=	"11" when vga_fb = '1' else 
				"10" when vga_ht = '1' else
				"00";
   vgab <=	"00";
   vgav <= vga_vsync;
   vgah <= vga_hsync;

   dram_match <= '1' when addr(21 downto 18) /= "1111" else '0';
   dram_cke <= '1';
   dram_clk <= c0;

   process(c0)
   begin
      if c0='1' and c0'event then
         if slowreset = '1' then
            dram_fsm <= dram_init;
            dram_cs_n <= '0';
            dram_ras_n <= '1';
            dram_cas_n <= '1';
            dram_we_n <= '1';
            dram_addr <= (others => '0');

            dram_udqm <= '1';
            dram_ldqm <= '1';
            dram_ba_1 <= '0';
            dram_ba_0 <= '0';

            cpuclk <= '0';
            cpureset <= '1';
            cpuresetlength <= 63;
				-- Select the drive type from jumpers
            if sw(2 downto 0) = "110" then
               have_rl <= 1;
               have_rk <= 0;
					have_rh <= 0;
            elsif sw(2 downto 0) = "101" then
               have_rl <= 0;
               have_rk <= 1;
					have_rh <= 0;
            elsif sw(2 downto 0) = "011" then
               have_rl <= 0;
               have_rk <= 0;
					have_rh <= 1;
            end if;
				if sw(3) = '1' then 
					have_kl11 <= 1;
				else
					have_kl11 <= 0;
            end if;
				if sw(4) = '1' then 
					have_xu <= 1;
				else
					have_xu <= 0;
            end if;
         else

            case dram_fsm is

               when dram_init =>
                  dram_cs_n <= '0';
                  dram_ras_n <= '1';
                  dram_cas_n <= '1';
                  dram_we_n <= '1';
                  dram_addr <= (others => '0');

                  dram_udqm <= '1';
                  dram_ldqm <= '1';
                  dram_ba_1 <= '0';
                  dram_ba_0 <= '0';

                  cpureset <= '1';
                  cpuresetlength <= 8;
                  dram_counter <= 32767;
                  dram_fsm <= dram_poweron;

               when dram_poweron =>
                  dram_cs_n <= '0';
                  dram_ras_n <= '1';
                  dram_cas_n <= '1';
                  dram_we_n <= '1';
                  dram_addr <= (others => '0');

                  dram_udqm <= '1';
                  dram_ldqm <= '1';
                  dram_ba_1 <= '0';
                  dram_ba_0 <= '0';

                  if dram_counter = 0 then
                     dram_fsm <= dram_pwron_pre;
                  else
                     dram_counter <= dram_counter - 1;
                  end if;

               when dram_pwron_pre =>
                  dram_cs_n <= '0';
                  dram_ras_n <= '0';
                  dram_cas_n <= '1';
                  dram_we_n <= '0';
                  dram_addr(10) <= '1';

                  dram_udqm <= '1';
                  dram_ldqm <= '1';
                  dram_ba_1 <= '0';
                  dram_ba_0 <= '0';
                  dram_addr(12) <= '0';
                  dram_addr(11) <= '0';
                  dram_addr(9 downto 0) <= (others => '0');

                  dram_wait <= 4;
                  dram_fsm <= dram_pwron_prew;

               when dram_pwron_prew =>
                  dram_cs_n <= '1';
                  if dram_wait = 0 then
                     dram_fsm <= dram_pwron_ref;
                     dram_counter <= 20;
                  else
                     dram_wait <= dram_wait - 1;
                  end if;

               when dram_pwron_ref =>
                  dram_cs_n <= '0';
                  dram_ras_n <= '0';
                  dram_cas_n <= '0';
                  dram_we_n <= '1';
                  dram_addr <= (others => '0');

                  dram_udqm <= '1';
                  dram_ldqm <= '1';
                  dram_ba_1 <= '0';
                  dram_ba_0 <= '0';

                  dram_wait <= 15;
                  dram_fsm <= dram_pwron_refw;

               when dram_pwron_refw =>
                  dram_cs_n <= '1';
                  if dram_wait = 0 then
                     if dram_counter = 0 then
                        dram_fsm <= dram_pwron_mrs;
                     else
                        dram_counter <= dram_counter - 1;
                        dram_fsm <= dram_pwron_ref;
                     end if;
                  else
                     dram_wait <= dram_wait - 1;
                  end if;

               when dram_pwron_mrs =>
                  dram_cs_n <= '0';
                  dram_ras_n <= '0';
                  dram_cas_n <= '0';
                  dram_we_n <= '0';

                  dram_addr(12 downto 7) <= (others => '0');
                  dram_addr(6 downto 4) <= "011";          -- cas length 3
                  dram_addr(3) <= '0';                     -- sequential
                  dram_addr(2 downto 0) <= "000";          -- length 0

                  dram_udqm <= '1';
                  dram_ldqm <= '1';
                  dram_ba_1 <= '0';
                  dram_ba_0 <= '0';

                  dram_wait <= 4;
                  dram_fsm <= dram_pwron_mrsw;

               when dram_pwron_mrsw =>
                  dram_cs_n <= '1';
                  if dram_wait = 0 then
                     dram_fsm <= dram_idle;
                  else
                     dram_wait <= dram_wait - 1;
                  end if;

               when dram_idle =>
                  dram_cs_n <= '1';
                  dram_ras_n <= '1';
                  dram_cas_n <= '1';
                  dram_we_n <= '1';
                  dram_addr(10) <= '0';

                  dram_udqm <= '1';
                  dram_ldqm <= '1';
                  dram_ba_1 <= '0';
                  dram_ba_0 <= '0';
                  dram_addr(12) <= '0';
                  dram_addr(11) <= '0';
                  dram_addr(9 downto 0) <= (others => '0');

                  dram_fsm <= dram_c1;

               when dram_c1 =>

               cpuclk <= '1';

                  if cpuresetlength = 0 then
                     cpureset <= '0';
                  else
                     cpuresetlength <= cpuresetlength - 1;
                  end if;
                  dram_fsm <= dram_c2;

               when dram_c2 =>
                  dram_dq <= (others => 'Z');
                  dram_fsm <= dram_c3;

               when dram_c3 =>
                  dram_fsm <= dram_c4;

               when dram_c4 =>
                  dram_fsm <= dram_c5;

               when dram_c5 =>
                  dram_fsm <= dram_c6;

               when dram_c6 =>
                  -- read, t1-t2
                  if ifetch = '1' then
                     addrq <= addr;
                  end if;

                  if dram_match = '1' and control_dati = '1' then
                     -- activate command
                     dram_cs_n <= '0';
                     dram_ras_n <= '0';
                     dram_cas_n <= '1';
                     dram_we_n <= '1';
                     dram_addr(12) <= '0';
                     dram_addr(11 downto 0) <= addr(20 downto 9);

                     dram_udqm <= '0';
                     dram_ldqm <= '0';
                     dram_ba_1 <= '0';
                     dram_ba_0 <= addr(21);
                  end if;

                  -- write, t1-t2
                  if dram_match = '1' and control_dato = '1' then
                     -- activate command
                     dram_cs_n <= '0';
                     dram_ras_n <= '0';
                     dram_cas_n <= '1';
                     dram_we_n <= '1';
                     dram_addr(12) <= '0';
                     dram_addr(11 downto 0) <= addr(20 downto 9);

                     dram_udqm <= '0';
                     dram_ldqm <= '0';
                     dram_ba_1 <= '0';
                     dram_ba_0 <= addr(21);
                  end if;

                  if dram_match = '0' or (control_dato = '0' and control_dati = '0') then
                     -- auto refresh command
                     dram_cs_n <= '0';
                     dram_ras_n <= '0';
                     dram_cas_n <= '0';
                     dram_we_n <= '1';
                  end if;

                  dram_fsm <= dram_c7;

               when dram_c7 =>
                  -- t2-t3 - set nop command
                  dram_cs_n <= '1';
                  dram_ras_n <= '1';
                  dram_cas_n <= '1';
                  dram_we_n <= '1';

                  dram_fsm <= dram_c8;

               when dram_c8 =>

                  -- read, t3-t4
                  if dram_match = '1' and control_dati = '1' then
                     -- reada command
                     dram_cs_n <= '0';
                     dram_ras_n <= '1';
                     dram_cas_n <= '0';
                     dram_we_n <= '1';
                     dram_addr(12) <= '0';
                     dram_addr(11) <= '0';
                     dram_addr(10) <= '1';
                     dram_addr(9) <= '1';
                     dram_addr(8) <= '0';
                     dram_addr(7 downto 0) <= addr(8 downto 1);

                     dram_udqm <= '0';
                     dram_ldqm <= '0';
                     dram_ba_1 <= '0';
                     dram_ba_0 <= addr(21);
                  end if;

                  -- write, t3-t4
                  if dram_match = '1' and control_dato = '1' then
                     -- writea command
                     dram_cs_n <= '0';
                     dram_ras_n <= '1';
                     dram_cas_n <= '0';
                     dram_we_n <= '0';
                     dram_addr(12) <= '0';
                     dram_addr(11) <= '0';
                     dram_addr(10) <= '1';
                     dram_addr(9) <= '1';
                     dram_addr(8) <= '0';
                     dram_addr(7 downto 0) <= addr(8 downto 1);
                     dram_udqm <= '0';
                     dram_ldqm <= '0';
                     if control_datob = '1' then
                        if addr(0) = '0' then
                           dram_udqm <= '1';
                        else
                           dram_ldqm <= '1';
                        end if;
                     end if;
                     dram_ba_1 <= '0';
                     dram_ba_0 <= addr(21);
                     dram_dq <= dato;
                  end if;

                  dram_fsm <= dram_c9;

               cpuclk <= '0';

               when dram_c9 =>
                  -- read/write, t4-t5 - set nop command and deselect
                  dram_cs_n <= '1';
                  dram_ras_n <= '1';
                  dram_cas_n <= '1';
                  dram_we_n <= '1';

                  dram_fsm <= dram_c10;

               when dram_c10 =>
                  dram_fsm <= dram_c11;

               when dram_c11 =>
                  dram_fsm <= dram_c12;

               when dram_c12 =>
                  dram_fsm <= dram_c13;

               when dram_c13 =>
                  -- read, t5-t6
                  if dram_match = '1' and control_dati = '1' then
                     dati <= dram_dq;
                  end if;
                  dram_fsm <= dram_c14;

               when dram_c14 =>
                  dram_fsm <= dram_c1;

               when others =>
                  null;

            end case;

         end if;
      end if;
   end process;

   process (c0)
   begin
      if c0='1' and c0'event then
         if reset = '1' then
            slowreset <= '1';
            slowresetdelay <= 4095;
         else
            if slowresetdelay = 0 then
               slowreset <= '0';
               vtreset <= '0';
            else
               slowreset <= '1';
               slowresetdelay <= slowresetdelay - 1;
            end if;
         end if;
      end if;
   end process;

end implementation;

