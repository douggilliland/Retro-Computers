library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity CharROM_ROM is
generic
	(
		addrbits : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clock : in std_logic;
	address : in std_logic_vector(addrbits-1 downto 0);
	q : out std_logic_vector(7 downto 0)
);
end CharROM_ROM;

architecture arch of CharROM_ROM is

type rom_type is array(natural range 0 to (2**(addrbits)-1)) of std_logic_vector(7 downto 0);

shared variable rom : rom_type :=
(
     0 => x"00",
     1 => x"00",
     2 => x"00",
     3 => x"00",
     4 => x"00",
     5 => x"00",
     6 => x"00",
     7 => x"00",
     8 => x"00",
     9 => x"00",
    10 => x"00",
    11 => x"00",
    12 => x"00",
    13 => x"00",
    14 => x"00",
    15 => x"00",
    16 => x"00",
    17 => x"00",
    18 => x"00",
    19 => x"00",
    20 => x"00",
    21 => x"00",
    22 => x"00",
    23 => x"00",
    24 => x"00",
    25 => x"00",
    26 => x"00",
    27 => x"00",
    28 => x"00",
    29 => x"00",
    30 => x"00",
    31 => x"00",
    32 => x"00",
    33 => x"00",
    34 => x"00",
    35 => x"00",
    36 => x"00",
    37 => x"00",
    38 => x"00",
    39 => x"00",
    40 => x"00",
    41 => x"00",
    42 => x"00",
    43 => x"00",
    44 => x"00",
    45 => x"00",
    46 => x"00",
    47 => x"00",
    48 => x"00",
    49 => x"00",
    50 => x"00",
    51 => x"00",
    52 => x"00",
    53 => x"00",
    54 => x"00",
    55 => x"00",
    56 => x"00",
    57 => x"00",
    58 => x"00",
    59 => x"00",
    60 => x"00",
    61 => x"00",
    62 => x"00",
    63 => x"00",
    64 => x"00",
    65 => x"00",
    66 => x"00",
    67 => x"00",
    68 => x"00",
    69 => x"00",
    70 => x"00",
    71 => x"00",
    72 => x"00",
    73 => x"00",
    74 => x"00",
    75 => x"00",
    76 => x"00",
    77 => x"00",
    78 => x"00",
    79 => x"00",
    80 => x"00",
    81 => x"00",
    82 => x"00",
    83 => x"00",
    84 => x"00",
    85 => x"00",
    86 => x"00",
    87 => x"00",
    88 => x"00",
    89 => x"00",
    90 => x"00",
    91 => x"00",
    92 => x"00",
    93 => x"00",
    94 => x"00",
    95 => x"00",
    96 => x"00",
    97 => x"00",
    98 => x"00",
    99 => x"00",
   100 => x"00",
   101 => x"00",
   102 => x"00",
   103 => x"00",
   104 => x"00",
   105 => x"00",
   106 => x"00",
   107 => x"00",
   108 => x"00",
   109 => x"00",
   110 => x"00",
   111 => x"00",
   112 => x"00",
   113 => x"00",
   114 => x"00",
   115 => x"00",
   116 => x"00",
   117 => x"00",
   118 => x"00",
   119 => x"00",
   120 => x"00",
   121 => x"00",
   122 => x"00",
   123 => x"00",
   124 => x"00",
   125 => x"00",
   126 => x"00",
   127 => x"00",
   128 => x"00",
   129 => x"00",
   130 => x"00",
   131 => x"00",
   132 => x"00",
   133 => x"00",
   134 => x"00",
   135 => x"00",
   136 => x"00",
   137 => x"00",
   138 => x"00",
   139 => x"00",
   140 => x"00",
   141 => x"00",
   142 => x"00",
   143 => x"00",
   144 => x"00",
   145 => x"00",
   146 => x"00",
   147 => x"00",
   148 => x"00",
   149 => x"00",
   150 => x"00",
   151 => x"00",
   152 => x"00",
   153 => x"00",
   154 => x"00",
   155 => x"00",
   156 => x"00",
   157 => x"00",
   158 => x"00",
   159 => x"00",
   160 => x"00",
   161 => x"00",
   162 => x"00",
   163 => x"00",
   164 => x"00",
   165 => x"00",
   166 => x"00",
   167 => x"00",
   168 => x"00",
   169 => x"00",
   170 => x"00",
   171 => x"00",
   172 => x"00",
   173 => x"00",
   174 => x"00",
   175 => x"00",
   176 => x"00",
   177 => x"00",
   178 => x"00",
   179 => x"00",
   180 => x"00",
   181 => x"00",
   182 => x"00",
   183 => x"00",
   184 => x"00",
   185 => x"00",
   186 => x"00",
   187 => x"00",
   188 => x"00",
   189 => x"00",
   190 => x"00",
   191 => x"00",
   192 => x"00",
   193 => x"00",
   194 => x"00",
   195 => x"00",
   196 => x"00",
   197 => x"00",
   198 => x"00",
   199 => x"00",
   200 => x"00",
   201 => x"00",
   202 => x"00",
   203 => x"00",
   204 => x"00",
   205 => x"00",
   206 => x"00",
   207 => x"00",
   208 => x"00",
   209 => x"00",
   210 => x"00",
   211 => x"00",
   212 => x"00",
   213 => x"00",
   214 => x"00",
   215 => x"00",
   216 => x"00",
   217 => x"00",
   218 => x"00",
   219 => x"00",
   220 => x"00",
   221 => x"00",
   222 => x"00",
   223 => x"00",
   224 => x"00",
   225 => x"00",
   226 => x"00",
   227 => x"00",
   228 => x"00",
   229 => x"00",
   230 => x"00",
   231 => x"00",
   232 => x"00",
   233 => x"00",
   234 => x"00",
   235 => x"00",
   236 => x"00",
   237 => x"00",
   238 => x"00",
   239 => x"00",
   240 => x"00",
   241 => x"00",
   242 => x"00",
   243 => x"00",
   244 => x"00",
   245 => x"00",
   246 => x"00",
   247 => x"00",
   248 => x"00",
   249 => x"00",
   250 => x"00",
   251 => x"00",
   252 => x"00",
   253 => x"00",
   254 => x"00",
   255 => x"00",
   256 => x"00",
   257 => x"00",
   258 => x"00",
   259 => x"00",
   260 => x"00",
   261 => x"00",
   262 => x"00",
   263 => x"00",
   264 => x"18",
   265 => x"18",
   266 => x"18",
   267 => x"18",
   268 => x"18",
   269 => x"00",
   270 => x"18",
   271 => x"00",
   272 => x"6c",
   273 => x"6c",
   274 => x"00",
   275 => x"00",
   276 => x"00",
   277 => x"00",
   278 => x"00",
   279 => x"00",
   280 => x"6c",
   281 => x"6c",
   282 => x"fe",
   283 => x"6c",
   284 => x"fe",
   285 => x"6c",
   286 => x"6c",
   287 => x"00",
   288 => x"18",
   289 => x"3e",
   290 => x"60",
   291 => x"3c",
   292 => x"06",
   293 => x"7c",
   294 => x"18",
   295 => x"00",
   296 => x"00",
   297 => x"66",
   298 => x"ac",
   299 => x"d8",
   300 => x"36",
   301 => x"6a",
   302 => x"cc",
   303 => x"00",
   304 => x"38",
   305 => x"6c",
   306 => x"68",
   307 => x"76",
   308 => x"dc",
   309 => x"ce",
   310 => x"7b",
   311 => x"00",
   312 => x"18",
   313 => x"18",
   314 => x"30",
   315 => x"00",
   316 => x"00",
   317 => x"00",
   318 => x"00",
   319 => x"00",
   320 => x"0c",
   321 => x"18",
   322 => x"30",
   323 => x"30",
   324 => x"30",
   325 => x"18",
   326 => x"0c",
   327 => x"00",
   328 => x"30",
   329 => x"18",
   330 => x"0c",
   331 => x"0c",
   332 => x"0c",
   333 => x"18",
   334 => x"30",
   335 => x"00",
   336 => x"00",
   337 => x"66",
   338 => x"3c",
   339 => x"ff",
   340 => x"3c",
   341 => x"66",
   342 => x"00",
   343 => x"00",
   344 => x"00",
   345 => x"18",
   346 => x"18",
   347 => x"7e",
   348 => x"18",
   349 => x"18",
   350 => x"00",
   351 => x"00",
   352 => x"00",
   353 => x"00",
   354 => x"00",
   355 => x"00",
   356 => x"00",
   357 => x"18",
   358 => x"18",
   359 => x"30",
   360 => x"00",
   361 => x"00",
   362 => x"00",
   363 => x"7e",
   364 => x"00",
   365 => x"00",
   366 => x"00",
   367 => x"00",
   368 => x"00",
   369 => x"00",
   370 => x"00",
   371 => x"00",
   372 => x"00",
   373 => x"18",
   374 => x"18",
   375 => x"00",
   376 => x"03",
   377 => x"06",
   378 => x"0c",
   379 => x"18",
   380 => x"30",
   381 => x"60",
   382 => x"c0",
   383 => x"00",
   384 => x"3c",
   385 => x"66",
   386 => x"6e",
   387 => x"7e",
   388 => x"76",
   389 => x"66",
   390 => x"3c",
   391 => x"00",
   392 => x"18",
   393 => x"38",
   394 => x"78",
   395 => x"18",
   396 => x"18",
   397 => x"18",
   398 => x"18",
   399 => x"00",
   400 => x"3c",
   401 => x"66",
   402 => x"06",
   403 => x"0c",
   404 => x"18",
   405 => x"30",
   406 => x"7e",
   407 => x"00",
   408 => x"3c",
   409 => x"66",
   410 => x"06",
   411 => x"1c",
   412 => x"06",
   413 => x"66",
   414 => x"3c",
   415 => x"00",
   416 => x"1c",
   417 => x"3c",
   418 => x"6c",
   419 => x"cc",
   420 => x"fe",
   421 => x"0c",
   422 => x"0c",
   423 => x"00",
   424 => x"7e",
   425 => x"60",
   426 => x"7c",
   427 => x"06",
   428 => x"06",
   429 => x"66",
   430 => x"3c",
   431 => x"00",
   432 => x"1c",
   433 => x"30",
   434 => x"60",
   435 => x"7c",
   436 => x"66",
   437 => x"66",
   438 => x"3c",
   439 => x"00",
   440 => x"7e",
   441 => x"06",
   442 => x"06",
   443 => x"0c",
   444 => x"18",
   445 => x"18",
   446 => x"18",
   447 => x"00",
   448 => x"3c",
   449 => x"66",
   450 => x"66",
   451 => x"3c",
   452 => x"66",
   453 => x"66",
   454 => x"3c",
   455 => x"00",
   456 => x"3c",
   457 => x"66",
   458 => x"66",
   459 => x"3e",
   460 => x"06",
   461 => x"0c",
   462 => x"38",
   463 => x"00",
   464 => x"00",
   465 => x"18",
   466 => x"18",
   467 => x"00",
   468 => x"00",
   469 => x"18",
   470 => x"18",
   471 => x"00",
   472 => x"00",
   473 => x"18",
   474 => x"18",
   475 => x"00",
   476 => x"00",
   477 => x"18",
   478 => x"18",
   479 => x"30",
   480 => x"00",
   481 => x"06",
   482 => x"18",
   483 => x"60",
   484 => x"18",
   485 => x"06",
   486 => x"00",
   487 => x"00",
   488 => x"00",
   489 => x"00",
   490 => x"7e",
   491 => x"00",
   492 => x"7e",
   493 => x"00",
   494 => x"00",
   495 => x"00",
   496 => x"00",
   497 => x"60",
   498 => x"18",
   499 => x"06",
   500 => x"18",
   501 => x"60",
   502 => x"00",
   503 => x"00",
   504 => x"3c",
   505 => x"66",
   506 => x"06",
   507 => x"0c",
   508 => x"18",
   509 => x"00",
   510 => x"18",
   511 => x"00",
   512 => x"7c",
   513 => x"c6",
   514 => x"de",
   515 => x"d6",
   516 => x"de",
   517 => x"c0",
   518 => x"78",
   519 => x"00",
   520 => x"3c",
   521 => x"66",
   522 => x"66",
   523 => x"7e",
   524 => x"66",
   525 => x"66",
   526 => x"66",
   527 => x"00",
   528 => x"7c",
   529 => x"66",
   530 => x"66",
   531 => x"7c",
   532 => x"66",
   533 => x"66",
   534 => x"7c",
   535 => x"00",
   536 => x"1e",
   537 => x"30",
   538 => x"60",
   539 => x"60",
   540 => x"60",
   541 => x"30",
   542 => x"1e",
   543 => x"00",
   544 => x"78",
   545 => x"6c",
   546 => x"66",
   547 => x"66",
   548 => x"66",
   549 => x"6c",
   550 => x"78",
   551 => x"00",
   552 => x"7e",
   553 => x"60",
   554 => x"60",
   555 => x"78",
   556 => x"60",
   557 => x"60",
   558 => x"7e",
   559 => x"00",
   560 => x"7e",
   561 => x"60",
   562 => x"60",
   563 => x"78",
   564 => x"60",
   565 => x"60",
   566 => x"60",
   567 => x"00",
   568 => x"3c",
   569 => x"66",
   570 => x"60",
   571 => x"6e",
   572 => x"66",
   573 => x"66",
   574 => x"3e",
   575 => x"00",
   576 => x"66",
   577 => x"66",
   578 => x"66",
   579 => x"7e",
   580 => x"66",
   581 => x"66",
   582 => x"66",
   583 => x"00",
   584 => x"3c",
   585 => x"18",
   586 => x"18",
   587 => x"18",
   588 => x"18",
   589 => x"18",
   590 => x"3c",
   591 => x"00",
   592 => x"06",
   593 => x"06",
   594 => x"06",
   595 => x"06",
   596 => x"06",
   597 => x"66",
   598 => x"3c",
   599 => x"00",
   600 => x"c6",
   601 => x"cc",
   602 => x"d8",
   603 => x"f0",
   604 => x"d8",
   605 => x"cc",
   606 => x"c6",
   607 => x"00",
   608 => x"60",
   609 => x"60",
   610 => x"60",
   611 => x"60",
   612 => x"60",
   613 => x"60",
   614 => x"7e",
   615 => x"00",
   616 => x"c6",
   617 => x"ee",
   618 => x"fe",
   619 => x"d6",
   620 => x"c6",
   621 => x"c6",
   622 => x"c6",
   623 => x"00",
   624 => x"c6",
   625 => x"e6",
   626 => x"f6",
   627 => x"de",
   628 => x"ce",
   629 => x"c6",
   630 => x"c6",
   631 => x"00",
   632 => x"3c",
   633 => x"66",
   634 => x"66",
   635 => x"66",
   636 => x"66",
   637 => x"66",
   638 => x"3c",
   639 => x"00",
   640 => x"7c",
   641 => x"66",
   642 => x"66",
   643 => x"7c",
   644 => x"60",
   645 => x"60",
   646 => x"60",
   647 => x"00",
   648 => x"78",
   649 => x"cc",
   650 => x"cc",
   651 => x"cc",
   652 => x"cc",
   653 => x"dc",
   654 => x"7e",
   655 => x"00",
   656 => x"7c",
   657 => x"66",
   658 => x"66",
   659 => x"7c",
   660 => x"6c",
   661 => x"66",
   662 => x"66",
   663 => x"00",
   664 => x"3c",
   665 => x"66",
   666 => x"70",
   667 => x"3c",
   668 => x"0e",
   669 => x"66",
   670 => x"3c",
   671 => x"00",
   672 => x"7e",
   673 => x"18",
   674 => x"18",
   675 => x"18",
   676 => x"18",
   677 => x"18",
   678 => x"18",
   679 => x"00",
   680 => x"66",
   681 => x"66",
   682 => x"66",
   683 => x"66",
   684 => x"66",
   685 => x"66",
   686 => x"3c",
   687 => x"00",
   688 => x"66",
   689 => x"66",
   690 => x"66",
   691 => x"66",
   692 => x"3c",
   693 => x"3c",
   694 => x"18",
   695 => x"00",
   696 => x"c6",
   697 => x"c6",
   698 => x"c6",
   699 => x"d6",
   700 => x"fe",
   701 => x"ee",
   702 => x"c6",
   703 => x"00",
   704 => x"c3",
   705 => x"66",
   706 => x"3c",
   707 => x"18",
   708 => x"3c",
   709 => x"66",
   710 => x"c3",
   711 => x"00",
   712 => x"c3",
   713 => x"66",
   714 => x"3c",
   715 => x"18",
   716 => x"18",
   717 => x"18",
   718 => x"18",
   719 => x"00",
   720 => x"fe",
   721 => x"0c",
   722 => x"18",
   723 => x"30",
   724 => x"60",
   725 => x"c0",
   726 => x"fe",
   727 => x"00",
   728 => x"3c",
   729 => x"30",
   730 => x"30",
   731 => x"30",
   732 => x"30",
   733 => x"30",
   734 => x"3c",
   735 => x"00",
   736 => x"c0",
   737 => x"60",
   738 => x"30",
   739 => x"18",
   740 => x"0c",
   741 => x"06",
   742 => x"03",
   743 => x"00",
   744 => x"3c",
   745 => x"0c",
   746 => x"0c",
   747 => x"0c",
   748 => x"0c",
   749 => x"0c",
   750 => x"3c",
   751 => x"00",
   752 => x"10",
   753 => x"38",
   754 => x"6c",
   755 => x"c6",
   756 => x"00",
   757 => x"00",
   758 => x"00",
   759 => x"00",
   760 => x"00",
   761 => x"00",
   762 => x"00",
   763 => x"00",
   764 => x"00",
   765 => x"00",
   766 => x"00",
   767 => x"fe",
   768 => x"18",
   769 => x"18",
   770 => x"0c",
   771 => x"00",
   772 => x"00",
   773 => x"00",
   774 => x"00",
   775 => x"00",
   776 => x"00",
   777 => x"00",
   778 => x"3c",
   779 => x"06",
   780 => x"3e",
   781 => x"66",
   782 => x"3e",
   783 => x"00",
   784 => x"60",
   785 => x"60",
   786 => x"7c",
   787 => x"66",
   788 => x"66",
   789 => x"66",
   790 => x"7c",
   791 => x"00",
   792 => x"00",
   793 => x"00",
   794 => x"3c",
   795 => x"60",
   796 => x"60",
   797 => x"60",
   798 => x"3c",
   799 => x"00",
   800 => x"06",
   801 => x"06",
   802 => x"3e",
   803 => x"66",
   804 => x"66",
   805 => x"66",
   806 => x"3e",
   807 => x"00",
   808 => x"00",
   809 => x"00",
   810 => x"3c",
   811 => x"66",
   812 => x"7e",
   813 => x"60",
   814 => x"3c",
   815 => x"00",
   816 => x"1c",
   817 => x"30",
   818 => x"7c",
   819 => x"30",
   820 => x"30",
   821 => x"30",
   822 => x"30",
   823 => x"00",
   824 => x"00",
   825 => x"00",
   826 => x"3e",
   827 => x"66",
   828 => x"66",
   829 => x"3e",
   830 => x"06",
   831 => x"3c",
   832 => x"60",
   833 => x"60",
   834 => x"7c",
   835 => x"66",
   836 => x"66",
   837 => x"66",
   838 => x"66",
   839 => x"00",
   840 => x"18",
   841 => x"00",
   842 => x"18",
   843 => x"18",
   844 => x"18",
   845 => x"18",
   846 => x"0c",
   847 => x"00",
   848 => x"0c",
   849 => x"00",
   850 => x"0c",
   851 => x"0c",
   852 => x"0c",
   853 => x"0c",
   854 => x"0c",
   855 => x"78",
   856 => x"60",
   857 => x"60",
   858 => x"66",
   859 => x"6c",
   860 => x"78",
   861 => x"6c",
   862 => x"66",
   863 => x"00",
   864 => x"18",
   865 => x"18",
   866 => x"18",
   867 => x"18",
   868 => x"18",
   869 => x"18",
   870 => x"0c",
   871 => x"00",
   872 => x"00",
   873 => x"00",
   874 => x"ec",
   875 => x"fe",
   876 => x"d6",
   877 => x"c6",
   878 => x"c6",
   879 => x"00",
   880 => x"00",
   881 => x"00",
   882 => x"7c",
   883 => x"66",
   884 => x"66",
   885 => x"66",
   886 => x"66",
   887 => x"00",
   888 => x"00",
   889 => x"00",
   890 => x"3c",
   891 => x"66",
   892 => x"66",
   893 => x"66",
   894 => x"3c",
   895 => x"00",
   896 => x"00",
   897 => x"00",
   898 => x"7c",
   899 => x"66",
   900 => x"66",
   901 => x"7c",
   902 => x"60",
   903 => x"60",
   904 => x"00",
   905 => x"00",
   906 => x"3e",
   907 => x"66",
   908 => x"66",
   909 => x"3e",
   910 => x"06",
   911 => x"06",
   912 => x"00",
   913 => x"00",
   914 => x"7c",
   915 => x"66",
   916 => x"60",
   917 => x"60",
   918 => x"60",
   919 => x"00",
   920 => x"00",
   921 => x"00",
   922 => x"3c",
   923 => x"60",
   924 => x"3c",
   925 => x"06",
   926 => x"7c",
   927 => x"00",
   928 => x"30",
   929 => x"30",
   930 => x"7c",
   931 => x"30",
   932 => x"30",
   933 => x"30",
   934 => x"1c",
   935 => x"00",
   936 => x"00",
   937 => x"00",
   938 => x"66",
   939 => x"66",
   940 => x"66",
   941 => x"66",
   942 => x"3e",
   943 => x"00",
   944 => x"00",
   945 => x"00",
   946 => x"66",
   947 => x"66",
   948 => x"66",
   949 => x"3c",
   950 => x"18",
   951 => x"00",
   952 => x"00",
   953 => x"00",
   954 => x"c6",
   955 => x"c6",
   956 => x"d6",
   957 => x"fe",
   958 => x"6c",
   959 => x"00",
   960 => x"00",
   961 => x"00",
   962 => x"c6",
   963 => x"6c",
   964 => x"38",
   965 => x"6c",
   966 => x"c6",
   967 => x"00",
   968 => x"00",
   969 => x"00",
   970 => x"66",
   971 => x"66",
   972 => x"66",
   973 => x"3c",
   974 => x"18",
   975 => x"30",
   976 => x"00",
   977 => x"00",
   978 => x"7e",
   979 => x"0c",
   980 => x"18",
   981 => x"30",
   982 => x"7e",
   983 => x"00",
   984 => x"0e",
   985 => x"18",
   986 => x"18",
   987 => x"70",
   988 => x"18",
   989 => x"18",
   990 => x"0e",
   991 => x"00",
   992 => x"18",
   993 => x"18",
   994 => x"18",
   995 => x"18",
   996 => x"18",
   997 => x"18",
   998 => x"18",
   999 => x"00",
  1000 => x"70",
  1001 => x"18",
  1002 => x"18",
  1003 => x"0e",
  1004 => x"18",
  1005 => x"18",
  1006 => x"70",
  1007 => x"00",
  1008 => x"72",
  1009 => x"9c",
  1010 => x"00",
  1011 => x"00",
  1012 => x"00",
  1013 => x"00",
  1014 => x"00",
  1015 => x"00",
  1016 => x"fe",
  1017 => x"fe",
  1018 => x"fe",
  1019 => x"fe",
  1020 => x"fe",
  1021 => x"fe",
  1022 => x"fe",
  1023 => x"00",
	others => x"00"
);

begin

process (clock)
begin
	if (clock'event and clock = '1') then
		q(7 downto 0) <= rom(to_integer(unsigned(address(addrbits-1 downto 0))));
	end if;
end process;

end arch;

