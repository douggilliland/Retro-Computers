library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SanityCheck_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end SanityCheck_ROM;

architecture arch of SanityCheck_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"00",
     2 => x"0f",
     3 => x"fe",
     4 => x"00",
     5 => x"00",
     6 => x"01",
     7 => x"00",
     8 => x"00",
     9 => x"00",
    10 => x"00",
    11 => x"00",
    12 => x"00",
    13 => x"00",
    14 => x"00",
    15 => x"00",
    16 => x"00",
    17 => x"00",
    18 => x"00",
    19 => x"00",
    20 => x"00",
    21 => x"00",
    22 => x"00",
    23 => x"00",
    24 => x"00",
    25 => x"00",
    26 => x"00",
    27 => x"00",
    28 => x"00",
    29 => x"00",
    30 => x"00",
    31 => x"00",
    32 => x"00",
    33 => x"00",
    34 => x"00",
    35 => x"00",
    36 => x"00",
    37 => x"00",
    38 => x"00",
    39 => x"00",
    40 => x"00",
    41 => x"00",
    42 => x"00",
    43 => x"00",
    44 => x"00",
    45 => x"00",
    46 => x"00",
    47 => x"00",
    48 => x"00",
    49 => x"00",
    50 => x"00",
    51 => x"00",
    52 => x"00",
    53 => x"00",
    54 => x"00",
    55 => x"00",
    56 => x"00",
    57 => x"00",
    58 => x"00",
    59 => x"00",
    60 => x"00",
    61 => x"00",
    62 => x"00",
    63 => x"00",
    64 => x"00",
    65 => x"00",
    66 => x"00",
    67 => x"00",
    68 => x"00",
    69 => x"00",
    70 => x"00",
    71 => x"00",
    72 => x"00",
    73 => x"00",
    74 => x"00",
    75 => x"00",
    76 => x"00",
    77 => x"00",
    78 => x"00",
    79 => x"00",
    80 => x"00",
    81 => x"00",
    82 => x"00",
    83 => x"00",
    84 => x"00",
    85 => x"00",
    86 => x"00",
    87 => x"00",
    88 => x"00",
    89 => x"00",
    90 => x"00",
    91 => x"00",
    92 => x"00",
    93 => x"00",
    94 => x"00",
    95 => x"00",
    96 => x"00",
    97 => x"00",
    98 => x"00",
    99 => x"00",
   100 => x"00",
   101 => x"00",
   102 => x"00",
   103 => x"00",
   104 => x"00",
   105 => x"00",
   106 => x"00",
   107 => x"00",
   108 => x"00",
   109 => x"00",
   110 => x"00",
   111 => x"00",
   112 => x"00",
   113 => x"00",
   114 => x"00",
   115 => x"00",
   116 => x"00",
   117 => x"00",
   118 => x"00",
   119 => x"00",
   120 => x"00",
   121 => x"00",
   122 => x"00",
   123 => x"00",
   124 => x"00",
   125 => x"00",
   126 => x"00",
   127 => x"00",
   128 => x"00",
   129 => x"00",
   130 => x"00",
   131 => x"00",
   132 => x"00",
   133 => x"00",
   134 => x"00",
   135 => x"00",
   136 => x"00",
   137 => x"00",
   138 => x"00",
   139 => x"00",
   140 => x"00",
   141 => x"00",
   142 => x"00",
   143 => x"00",
   144 => x"00",
   145 => x"00",
   146 => x"00",
   147 => x"00",
   148 => x"00",
   149 => x"00",
   150 => x"00",
   151 => x"00",
   152 => x"00",
   153 => x"00",
   154 => x"00",
   155 => x"00",
   156 => x"00",
   157 => x"00",
   158 => x"00",
   159 => x"00",
   160 => x"00",
   161 => x"00",
   162 => x"00",
   163 => x"00",
   164 => x"00",
   165 => x"00",
   166 => x"00",
   167 => x"00",
   168 => x"00",
   169 => x"00",
   170 => x"00",
   171 => x"00",
   172 => x"00",
   173 => x"00",
   174 => x"00",
   175 => x"00",
   176 => x"00",
   177 => x"00",
   178 => x"00",
   179 => x"00",
   180 => x"00",
   181 => x"00",
   182 => x"00",
   183 => x"00",
   184 => x"00",
   185 => x"00",
   186 => x"00",
   187 => x"00",
   188 => x"00",
   189 => x"00",
   190 => x"00",
   191 => x"00",
   192 => x"00",
   193 => x"00",
   194 => x"00",
   195 => x"00",
   196 => x"00",
   197 => x"00",
   198 => x"00",
   199 => x"00",
   200 => x"00",
   201 => x"00",
   202 => x"00",
   203 => x"00",
   204 => x"00",
   205 => x"00",
   206 => x"00",
   207 => x"00",
   208 => x"00",
   209 => x"00",
   210 => x"00",
   211 => x"00",
   212 => x"00",
   213 => x"00",
   214 => x"00",
   215 => x"00",
   216 => x"00",
   217 => x"00",
   218 => x"00",
   219 => x"00",
   220 => x"00",
   221 => x"00",
   222 => x"00",
   223 => x"00",
   224 => x"00",
   225 => x"00",
   226 => x"00",
   227 => x"00",
   228 => x"00",
   229 => x"00",
   230 => x"00",
   231 => x"00",
   232 => x"00",
   233 => x"00",
   234 => x"00",
   235 => x"00",
   236 => x"00",
   237 => x"00",
   238 => x"00",
   239 => x"00",
   240 => x"00",
   241 => x"00",
   242 => x"00",
   243 => x"00",
   244 => x"00",
   245 => x"00",
   246 => x"00",
   247 => x"00",
   248 => x"00",
   249 => x"00",
   250 => x"00",
   251 => x"00",
   252 => x"00",
   253 => x"00",
   254 => x"00",
   255 => x"00",
   256 => x"4f",
   257 => x"f9",
   258 => x"00",
   259 => x"00",
   260 => x"0f",
   261 => x"fe",
   262 => x"41",
   263 => x"f9",
   264 => x"00",
   265 => x"00",
   266 => x"0a",
   267 => x"e8",
   268 => x"20",
   269 => x"3c",
   270 => x"00",
   271 => x"00",
   272 => x"0a",
   273 => x"e8",
   274 => x"b1",
   275 => x"c0",
   276 => x"6c",
   277 => x"04",
   278 => x"42",
   279 => x"98",
   280 => x"60",
   281 => x"f8",
   282 => x"41",
   283 => x"fa",
   284 => x"00",
   285 => x"4e",
   286 => x"21",
   287 => x"c8",
   288 => x"00",
   289 => x"64",
   290 => x"41",
   291 => x"fa",
   292 => x"00",
   293 => x"54",
   294 => x"21",
   295 => x"c8",
   296 => x"00",
   297 => x"68",
   298 => x"41",
   299 => x"fa",
   300 => x"00",
   301 => x"5a",
   302 => x"21",
   303 => x"c8",
   304 => x"00",
   305 => x"6c",
   306 => x"41",
   307 => x"fa",
   308 => x"00",
   309 => x"60",
   310 => x"21",
   311 => x"c8",
   312 => x"00",
   313 => x"70",
   314 => x"41",
   315 => x"fa",
   316 => x"00",
   317 => x"66",
   318 => x"21",
   319 => x"c8",
   320 => x"00",
   321 => x"74",
   322 => x"41",
   323 => x"fa",
   324 => x"00",
   325 => x"6c",
   326 => x"21",
   327 => x"c8",
   328 => x"00",
   329 => x"78",
   330 => x"41",
   331 => x"fa",
   332 => x"00",
   333 => x"72",
   334 => x"21",
   335 => x"c8",
   336 => x"00",
   337 => x"7c",
   338 => x"48",
   339 => x"78",
   340 => x"00",
   341 => x"01",
   342 => x"48",
   343 => x"7a",
   344 => x"00",
   345 => x"0a",
   346 => x"4e",
   347 => x"b9",
   348 => x"00",
   349 => x"00",
   350 => x"01",
   351 => x"fc",
   352 => x"60",
   353 => x"fe",
   354 => x"42",
   355 => x"6f",
   356 => x"6f",
   357 => x"74",
   358 => x"72",
   359 => x"6f",
   360 => x"6d",
   361 => x"00",
   362 => x"48",
   363 => x"e7",
   364 => x"ff",
   365 => x"fe",
   366 => x"48",
   367 => x"7a",
   368 => x"00",
   369 => x"5c",
   370 => x"2f",
   371 => x"3a",
   372 => x"00",
   373 => x"60",
   374 => x"4e",
   375 => x"75",
   376 => x"48",
   377 => x"e7",
   378 => x"ff",
   379 => x"fe",
   380 => x"48",
   381 => x"7a",
   382 => x"00",
   383 => x"4e",
   384 => x"2f",
   385 => x"3a",
   386 => x"00",
   387 => x"56",
   388 => x"4e",
   389 => x"75",
   390 => x"48",
   391 => x"e7",
   392 => x"ff",
   393 => x"fe",
   394 => x"48",
   395 => x"7a",
   396 => x"00",
   397 => x"40",
   398 => x"2f",
   399 => x"3a",
   400 => x"00",
   401 => x"4c",
   402 => x"4e",
   403 => x"75",
   404 => x"48",
   405 => x"e7",
   406 => x"ff",
   407 => x"fe",
   408 => x"48",
   409 => x"7a",
   410 => x"00",
   411 => x"32",
   412 => x"2f",
   413 => x"3a",
   414 => x"00",
   415 => x"42",
   416 => x"4e",
   417 => x"75",
   418 => x"48",
   419 => x"e7",
   420 => x"ff",
   421 => x"fe",
   422 => x"48",
   423 => x"7a",
   424 => x"00",
   425 => x"24",
   426 => x"2f",
   427 => x"3a",
   428 => x"00",
   429 => x"38",
   430 => x"4e",
   431 => x"75",
   432 => x"48",
   433 => x"e7",
   434 => x"ff",
   435 => x"fe",
   436 => x"48",
   437 => x"7a",
   438 => x"00",
   439 => x"16",
   440 => x"2f",
   441 => x"3a",
   442 => x"00",
   443 => x"2e",
   444 => x"4e",
   445 => x"75",
   446 => x"48",
   447 => x"e7",
   448 => x"ff",
   449 => x"fe",
   450 => x"48",
   451 => x"7a",
   452 => x"00",
   453 => x"08",
   454 => x"2f",
   455 => x"3a",
   456 => x"00",
   457 => x"24",
   458 => x"4e",
   459 => x"75",
   460 => x"4c",
   461 => x"df",
   462 => x"7f",
   463 => x"ff",
   464 => x"4e",
   465 => x"73",
   466 => x"4e",
   467 => x"75",
   468 => x"00",
   469 => x"00",
   470 => x"01",
   471 => x"d2",
   472 => x"00",
   473 => x"00",
   474 => x"01",
   475 => x"d2",
   476 => x"00",
   477 => x"00",
   478 => x"01",
   479 => x"d2",
   480 => x"00",
   481 => x"00",
   482 => x"01",
   483 => x"d2",
   484 => x"00",
   485 => x"00",
   486 => x"01",
   487 => x"d2",
   488 => x"00",
   489 => x"00",
   490 => x"01",
   491 => x"d2",
   492 => x"00",
   493 => x"00",
   494 => x"01",
   495 => x"d2",
   496 => x"46",
   497 => x"fc",
   498 => x"20",
   499 => x"00",
   500 => x"4e",
   501 => x"75",
   502 => x"46",
   503 => x"fc",
   504 => x"27",
   505 => x"00",
   506 => x"4e",
   507 => x"75",
   508 => x"4e",
   509 => x"56",
   510 => x"00",
   511 => x"00",
   512 => x"2f",
   513 => x"0a",
   514 => x"2f",
   515 => x"02",
   516 => x"32",
   517 => x"39",
   518 => x"81",
   519 => x"00",
   520 => x"00",
   521 => x"2a",
   522 => x"02",
   523 => x"81",
   524 => x"00",
   525 => x"00",
   526 => x"ff",
   527 => x"ff",
   528 => x"24",
   529 => x"01",
   530 => x"e5",
   531 => x"8a",
   532 => x"20",
   533 => x"01",
   534 => x"ef",
   535 => x"88",
   536 => x"90",
   537 => x"82",
   538 => x"d2",
   539 => x"80",
   540 => x"e7",
   541 => x"89",
   542 => x"24",
   543 => x"01",
   544 => x"4c",
   545 => x"3c",
   546 => x"2c",
   547 => x"00",
   548 => x"38",
   549 => x"e3",
   550 => x"8e",
   551 => x"39",
   552 => x"e0",
   553 => x"80",
   554 => x"d2",
   555 => x"81",
   556 => x"93",
   557 => x"81",
   558 => x"90",
   559 => x"81",
   560 => x"33",
   561 => x"c0",
   562 => x"81",
   563 => x"00",
   564 => x"00",
   565 => x"02",
   566 => x"48",
   567 => x"79",
   568 => x"00",
   569 => x"00",
   570 => x"0a",
   571 => x"a0",
   572 => x"45",
   573 => x"f9",
   574 => x"00",
   575 => x"00",
   576 => x"08",
   577 => x"06",
   578 => x"4e",
   579 => x"92",
   580 => x"2f",
   581 => x"3c",
   582 => x"00",
   583 => x"01",
   584 => x"00",
   585 => x"00",
   586 => x"4e",
   587 => x"b9",
   588 => x"00",
   589 => x"00",
   590 => x"06",
   591 => x"7a",
   592 => x"50",
   593 => x"8f",
   594 => x"4a",
   595 => x"80",
   596 => x"67",
   597 => x"08",
   598 => x"48",
   599 => x"79",
   600 => x"00",
   601 => x"00",
   602 => x"0a",
   603 => x"bd",
   604 => x"60",
   605 => x"06",
   606 => x"48",
   607 => x"79",
   608 => x"00",
   609 => x"00",
   610 => x"0a",
   611 => x"d2",
   612 => x"4e",
   613 => x"92",
   614 => x"58",
   615 => x"8f",
   616 => x"42",
   617 => x"80",
   618 => x"24",
   619 => x"2e",
   620 => x"ff",
   621 => x"f8",
   622 => x"24",
   623 => x"6e",
   624 => x"ff",
   625 => x"fc",
   626 => x"4e",
   627 => x"5e",
   628 => x"4e",
   629 => x"75",
   630 => x"00",
   631 => x"00",
   632 => x"4e",
   633 => x"56",
   634 => x"00",
   635 => x"00",
   636 => x"48",
   637 => x"e7",
   638 => x"38",
   639 => x"20",
   640 => x"24",
   641 => x"2e",
   642 => x"00",
   643 => x"08",
   644 => x"67",
   645 => x"3a",
   646 => x"76",
   647 => x"08",
   648 => x"42",
   649 => x"80",
   650 => x"45",
   651 => x"f9",
   652 => x"00",
   653 => x"00",
   654 => x"07",
   655 => x"e8",
   656 => x"22",
   657 => x"02",
   658 => x"78",
   659 => x"1c",
   660 => x"e8",
   661 => x"a9",
   662 => x"20",
   663 => x"41",
   664 => x"e9",
   665 => x"8a",
   666 => x"4a",
   667 => x"81",
   668 => x"67",
   669 => x"0c",
   670 => x"70",
   671 => x"09",
   672 => x"b0",
   673 => x"81",
   674 => x"6c",
   675 => x"0a",
   676 => x"41",
   677 => x"e8",
   678 => x"00",
   679 => x"37",
   680 => x"60",
   681 => x"08",
   682 => x"4a",
   683 => x"80",
   684 => x"67",
   685 => x"0c",
   686 => x"41",
   687 => x"e8",
   688 => x"00",
   689 => x"30",
   690 => x"2f",
   691 => x"08",
   692 => x"4e",
   693 => x"92",
   694 => x"58",
   695 => x"8f",
   696 => x"70",
   697 => x"01",
   698 => x"53",
   699 => x"83",
   700 => x"66",
   701 => x"d2",
   702 => x"60",
   703 => x"0c",
   704 => x"48",
   705 => x"78",
   706 => x"00",
   707 => x"30",
   708 => x"4e",
   709 => x"b9",
   710 => x"00",
   711 => x"00",
   712 => x"07",
   713 => x"e8",
   714 => x"58",
   715 => x"8f",
   716 => x"48",
   717 => x"78",
   718 => x"00",
   719 => x"0a",
   720 => x"4e",
   721 => x"b9",
   722 => x"00",
   723 => x"00",
   724 => x"07",
   725 => x"e8",
   726 => x"42",
   727 => x"80",
   728 => x"4c",
   729 => x"ee",
   730 => x"04",
   731 => x"1c",
   732 => x"ff",
   733 => x"f0",
   734 => x"4e",
   735 => x"5e",
   736 => x"4e",
   737 => x"75",
   738 => x"4e",
   739 => x"56",
   740 => x"00",
   741 => x"00",
   742 => x"20",
   743 => x"6e",
   744 => x"00",
   745 => x"08",
   746 => x"20",
   747 => x"28",
   748 => x"40",
   749 => x"00",
   750 => x"20",
   751 => x"30",
   752 => x"01",
   753 => x"70",
   754 => x"00",
   755 => x"01",
   756 => x"00",
   757 => x"04",
   758 => x"20",
   759 => x"30",
   760 => x"01",
   761 => x"70",
   762 => x"00",
   763 => x"00",
   764 => x"80",
   765 => x"00",
   766 => x"20",
   767 => x"30",
   768 => x"01",
   769 => x"70",
   770 => x"00",
   771 => x"00",
   772 => x"c0",
   773 => x"0c",
   774 => x"20",
   775 => x"30",
   776 => x"01",
   777 => x"70",
   778 => x"00",
   779 => x"00",
   780 => x"c0",
   781 => x"04",
   782 => x"20",
   783 => x"30",
   784 => x"01",
   785 => x"70",
   786 => x"00",
   787 => x"00",
   788 => x"80",
   789 => x"0c",
   790 => x"20",
   791 => x"30",
   792 => x"01",
   793 => x"70",
   794 => x"00",
   795 => x"01",
   796 => x"00",
   797 => x"00",
   798 => x"20",
   799 => x"28",
   800 => x"40",
   801 => x"08",
   802 => x"4e",
   803 => x"5e",
   804 => x"4e",
   805 => x"75",
   806 => x"4e",
   807 => x"56",
   808 => x"00",
   809 => x"00",
   810 => x"48",
   811 => x"e7",
   812 => x"38",
   813 => x"20",
   814 => x"24",
   815 => x"6e",
   816 => x"00",
   817 => x"08",
   818 => x"22",
   819 => x"2e",
   820 => x"00",
   821 => x"0c",
   822 => x"20",
   823 => x"2e",
   824 => x"00",
   825 => x"10",
   826 => x"26",
   827 => x"01",
   828 => x"48",
   829 => x"43",
   830 => x"42",
   831 => x"43",
   832 => x"24",
   833 => x"00",
   834 => x"42",
   835 => x"42",
   836 => x"48",
   837 => x"42",
   838 => x"84",
   839 => x"83",
   840 => x"24",
   841 => x"81",
   842 => x"25",
   843 => x"40",
   844 => x"00",
   845 => x"04",
   846 => x"26",
   847 => x"2a",
   848 => x"00",
   849 => x"02",
   850 => x"b4",
   851 => x"83",
   852 => x"67",
   853 => x"18",
   854 => x"48",
   855 => x"79",
   856 => x"00",
   857 => x"00",
   858 => x"08",
   859 => x"32",
   860 => x"4e",
   861 => x"b9",
   862 => x"00",
   863 => x"00",
   864 => x"08",
   865 => x"06",
   866 => x"2f",
   867 => x"03",
   868 => x"4e",
   869 => x"ba",
   870 => x"ff",
   871 => x"12",
   872 => x"b5",
   873 => x"83",
   874 => x"50",
   875 => x"8f",
   876 => x"60",
   877 => x"02",
   878 => x"42",
   879 => x"83",
   880 => x"48",
   881 => x"6a",
   882 => x"00",
   883 => x"08",
   884 => x"4e",
   885 => x"ba",
   886 => x"ff",
   887 => x"6c",
   888 => x"28",
   889 => x"2a",
   890 => x"00",
   891 => x"02",
   892 => x"58",
   893 => x"8f",
   894 => x"b4",
   895 => x"84",
   896 => x"67",
   897 => x"18",
   898 => x"48",
   899 => x"79",
   900 => x"00",
   901 => x"00",
   902 => x"08",
   903 => x"59",
   904 => x"4e",
   905 => x"b9",
   906 => x"00",
   907 => x"00",
   908 => x"08",
   909 => x"06",
   910 => x"2f",
   911 => x"04",
   912 => x"4e",
   913 => x"ba",
   914 => x"fe",
   915 => x"e6",
   916 => x"b9",
   917 => x"82",
   918 => x"86",
   919 => x"82",
   920 => x"50",
   921 => x"8f",
   922 => x"20",
   923 => x"03",
   924 => x"4c",
   925 => x"ee",
   926 => x"04",
   927 => x"1c",
   928 => x"ff",
   929 => x"f0",
   930 => x"4e",
   931 => x"5e",
   932 => x"4e",
   933 => x"75",
   934 => x"4e",
   935 => x"56",
   936 => x"00",
   937 => x"00",
   938 => x"48",
   939 => x"e7",
   940 => x"3f",
   941 => x"20",
   942 => x"24",
   943 => x"6e",
   944 => x"00",
   945 => x"08",
   946 => x"2a",
   947 => x"2e",
   948 => x"00",
   949 => x"0c",
   950 => x"20",
   951 => x"2e",
   952 => x"00",
   953 => x"10",
   954 => x"3e",
   955 => x"00",
   956 => x"42",
   957 => x"83",
   958 => x"36",
   959 => x"00",
   960 => x"28",
   961 => x"05",
   962 => x"42",
   963 => x"44",
   964 => x"88",
   965 => x"83",
   966 => x"48",
   967 => x"43",
   968 => x"42",
   969 => x"43",
   970 => x"86",
   971 => x"45",
   972 => x"24",
   973 => x"85",
   974 => x"34",
   975 => x"80",
   976 => x"24",
   977 => x"12",
   978 => x"b6",
   979 => x"82",
   980 => x"67",
   981 => x"18",
   982 => x"48",
   983 => x"79",
   984 => x"00",
   985 => x"00",
   986 => x"08",
   987 => x"80",
   988 => x"4e",
   989 => x"b9",
   990 => x"00",
   991 => x"00",
   992 => x"08",
   993 => x"06",
   994 => x"2f",
   995 => x"02",
   996 => x"4e",
   997 => x"ba",
   998 => x"fe",
   999 => x"92",
  1000 => x"b7",
  1001 => x"82",
  1002 => x"50",
  1003 => x"8f",
  1004 => x"60",
  1005 => x"02",
  1006 => x"42",
  1007 => x"82",
  1008 => x"2f",
  1009 => x"0a",
  1010 => x"4e",
  1011 => x"ba",
  1012 => x"fe",
  1013 => x"ee",
  1014 => x"2c",
  1015 => x"12",
  1016 => x"58",
  1017 => x"8f",
  1018 => x"b6",
  1019 => x"86",
  1020 => x"67",
  1021 => x"18",
  1022 => x"48",
  1023 => x"79",
  1024 => x"00",
  1025 => x"00",
  1026 => x"08",
  1027 => x"a4",
  1028 => x"4e",
  1029 => x"b9",
  1030 => x"00",
  1031 => x"00",
  1032 => x"08",
  1033 => x"06",
  1034 => x"2f",
  1035 => x"06",
  1036 => x"4e",
  1037 => x"ba",
  1038 => x"fe",
  1039 => x"6a",
  1040 => x"bd",
  1041 => x"83",
  1042 => x"84",
  1043 => x"83",
  1044 => x"50",
  1045 => x"8f",
  1046 => x"25",
  1047 => x"45",
  1048 => x"00",
  1049 => x"04",
  1050 => x"35",
  1051 => x"47",
  1052 => x"00",
  1053 => x"06",
  1054 => x"26",
  1055 => x"2a",
  1056 => x"00",
  1057 => x"04",
  1058 => x"b8",
  1059 => x"83",
  1060 => x"67",
  1061 => x"18",
  1062 => x"48",
  1063 => x"79",
  1064 => x"00",
  1065 => x"00",
  1066 => x"08",
  1067 => x"c8",
  1068 => x"4e",
  1069 => x"b9",
  1070 => x"00",
  1071 => x"00",
  1072 => x"08",
  1073 => x"06",
  1074 => x"2f",
  1075 => x"03",
  1076 => x"4e",
  1077 => x"ba",
  1078 => x"fe",
  1079 => x"42",
  1080 => x"b9",
  1081 => x"83",
  1082 => x"84",
  1083 => x"83",
  1084 => x"50",
  1085 => x"8f",
  1086 => x"48",
  1087 => x"6a",
  1088 => x"00",
  1089 => x"04",
  1090 => x"4e",
  1091 => x"ba",
  1092 => x"fe",
  1093 => x"9e",
  1094 => x"26",
  1095 => x"2a",
  1096 => x"00",
  1097 => x"04",
  1098 => x"58",
  1099 => x"8f",
  1100 => x"b8",
  1101 => x"83",
  1102 => x"67",
  1103 => x"18",
  1104 => x"48",
  1105 => x"79",
  1106 => x"00",
  1107 => x"00",
  1108 => x"08",
  1109 => x"ec",
  1110 => x"4e",
  1111 => x"b9",
  1112 => x"00",
  1113 => x"00",
  1114 => x"08",
  1115 => x"06",
  1116 => x"2f",
  1117 => x"03",
  1118 => x"4e",
  1119 => x"ba",
  1120 => x"fe",
  1121 => x"18",
  1122 => x"b7",
  1123 => x"84",
  1124 => x"84",
  1125 => x"84",
  1126 => x"50",
  1127 => x"8f",
  1128 => x"20",
  1129 => x"02",
  1130 => x"4c",
  1131 => x"ee",
  1132 => x"04",
  1133 => x"fc",
  1134 => x"ff",
  1135 => x"e4",
  1136 => x"4e",
  1137 => x"5e",
  1138 => x"4e",
  1139 => x"75",
  1140 => x"4e",
  1141 => x"56",
  1142 => x"00",
  1143 => x"00",
  1144 => x"48",
  1145 => x"e7",
  1146 => x"3f",
  1147 => x"3c",
  1148 => x"24",
  1149 => x"6e",
  1150 => x"00",
  1151 => x"08",
  1152 => x"26",
  1153 => x"2e",
  1154 => x"00",
  1155 => x"0c",
  1156 => x"20",
  1157 => x"2e",
  1158 => x"00",
  1159 => x"10",
  1160 => x"42",
  1161 => x"84",
  1162 => x"18",
  1163 => x"00",
  1164 => x"72",
  1165 => x"ff",
  1166 => x"46",
  1167 => x"01",
  1168 => x"c2",
  1169 => x"83",
  1170 => x"82",
  1171 => x"84",
  1172 => x"28",
  1173 => x"41",
  1174 => x"2e",
  1175 => x"04",
  1176 => x"e1",
  1177 => x"8f",
  1178 => x"22",
  1179 => x"03",
  1180 => x"02",
  1181 => x"41",
  1182 => x"00",
  1183 => x"ff",
  1184 => x"8e",
  1185 => x"81",
  1186 => x"2c",
  1187 => x"04",
  1188 => x"48",
  1189 => x"46",
  1190 => x"42",
  1191 => x"46",
  1192 => x"22",
  1193 => x"03",
  1194 => x"02",
  1195 => x"81",
  1196 => x"ff",
  1197 => x"00",
  1198 => x"ff",
  1199 => x"ff",
  1200 => x"8c",
  1201 => x"81",
  1202 => x"2a",
  1203 => x"04",
  1204 => x"72",
  1205 => x"18",
  1206 => x"e3",
  1207 => x"ad",
  1208 => x"22",
  1209 => x"03",
  1210 => x"02",
  1211 => x"81",
  1212 => x"00",
  1213 => x"ff",
  1214 => x"ff",
  1215 => x"ff",
  1216 => x"8a",
  1217 => x"81",
  1218 => x"24",
  1219 => x"83",
  1220 => x"15",
  1221 => x"40",
  1222 => x"00",
  1223 => x"03",
  1224 => x"25",
  1225 => x"43",
  1226 => x"00",
  1227 => x"04",
  1228 => x"15",
  1229 => x"40",
  1230 => x"00",
  1231 => x"06",
  1232 => x"25",
  1233 => x"43",
  1234 => x"00",
  1235 => x"08",
  1236 => x"15",
  1237 => x"40",
  1238 => x"00",
  1239 => x"09",
  1240 => x"25",
  1241 => x"43",
  1242 => x"00",
  1243 => x"0c",
  1244 => x"15",
  1245 => x"40",
  1246 => x"00",
  1247 => x"0c",
  1248 => x"24",
  1249 => x"12",
  1250 => x"b9",
  1251 => x"c2",
  1252 => x"67",
  1253 => x"26",
  1254 => x"48",
  1255 => x"79",
  1256 => x"00",
  1257 => x"00",
  1258 => x"09",
  1259 => x"10",
  1260 => x"4e",
  1261 => x"b9",
  1262 => x"00",
  1263 => x"00",
  1264 => x"08",
  1265 => x"06",
  1266 => x"2f",
  1267 => x"02",
  1268 => x"47",
  1269 => x"fa",
  1270 => x"fd",
  1271 => x"82",
  1272 => x"4e",
  1273 => x"93",
  1274 => x"2f",
  1275 => x"03",
  1276 => x"4e",
  1277 => x"93",
  1278 => x"2f",
  1279 => x"04",
  1280 => x"4e",
  1281 => x"93",
  1282 => x"20",
  1283 => x"0c",
  1284 => x"b1",
  1285 => x"82",
  1286 => x"4f",
  1287 => x"ef",
  1288 => x"00",
  1289 => x"10",
  1290 => x"60",
  1291 => x"02",
  1292 => x"42",
  1293 => x"82",
  1294 => x"47",
  1295 => x"ea",
  1296 => x"00",
  1297 => x"08",
  1298 => x"2f",
  1299 => x"0b",
  1300 => x"4e",
  1301 => x"ba",
  1302 => x"fd",
  1303 => x"cc",
  1304 => x"2a",
  1305 => x"52",
  1306 => x"58",
  1307 => x"8f",
  1308 => x"b9",
  1309 => x"cd",
  1310 => x"67",
  1311 => x"2a",
  1312 => x"48",
  1313 => x"79",
  1314 => x"00",
  1315 => x"00",
  1316 => x"09",
  1317 => x"33",
  1318 => x"4e",
  1319 => x"b9",
  1320 => x"00",
  1321 => x"00",
  1322 => x"08",
  1323 => x"06",
  1324 => x"2f",
  1325 => x"0d",
  1326 => x"4e",
  1327 => x"ba",
  1328 => x"fd",
  1329 => x"48",
  1330 => x"2f",
  1331 => x"03",
  1332 => x"4e",
  1333 => x"ba",
  1334 => x"fd",
  1335 => x"42",
  1336 => x"2f",
  1337 => x"04",
  1338 => x"4e",
  1339 => x"ba",
  1340 => x"fd",
  1341 => x"3c",
  1342 => x"20",
  1343 => x"0c",
  1344 => x"22",
  1345 => x"0d",
  1346 => x"b3",
  1347 => x"80",
  1348 => x"84",
  1349 => x"80",
  1350 => x"4f",
  1351 => x"ef",
  1352 => x"00",
  1353 => x"10",
  1354 => x"28",
  1355 => x"6a",
  1356 => x"00",
  1357 => x"04",
  1358 => x"be",
  1359 => x"8c",
  1360 => x"67",
  1361 => x"26",
  1362 => x"48",
  1363 => x"79",
  1364 => x"00",
  1365 => x"00",
  1366 => x"09",
  1367 => x"56",
  1368 => x"4e",
  1369 => x"b9",
  1370 => x"00",
  1371 => x"00",
  1372 => x"08",
  1373 => x"06",
  1374 => x"2f",
  1375 => x"0c",
  1376 => x"4b",
  1377 => x"fa",
  1378 => x"fd",
  1379 => x"16",
  1380 => x"4e",
  1381 => x"95",
  1382 => x"2f",
  1383 => x"03",
  1384 => x"4e",
  1385 => x"95",
  1386 => x"2f",
  1387 => x"04",
  1388 => x"4e",
  1389 => x"95",
  1390 => x"20",
  1391 => x"0c",
  1392 => x"bf",
  1393 => x"80",
  1394 => x"84",
  1395 => x"80",
  1396 => x"4f",
  1397 => x"ef",
  1398 => x"00",
  1399 => x"10",
  1400 => x"2f",
  1401 => x"0b",
  1402 => x"4e",
  1403 => x"ba",
  1404 => x"fd",
  1405 => x"66",
  1406 => x"28",
  1407 => x"6a",
  1408 => x"00",
  1409 => x"04",
  1410 => x"58",
  1411 => x"8f",
  1412 => x"be",
  1413 => x"8c",
  1414 => x"67",
  1415 => x"26",
  1416 => x"48",
  1417 => x"79",
  1418 => x"00",
  1419 => x"00",
  1420 => x"09",
  1421 => x"79",
  1422 => x"4e",
  1423 => x"b9",
  1424 => x"00",
  1425 => x"00",
  1426 => x"08",
  1427 => x"06",
  1428 => x"2f",
  1429 => x"0c",
  1430 => x"4b",
  1431 => x"fa",
  1432 => x"fc",
  1433 => x"e0",
  1434 => x"4e",
  1435 => x"95",
  1436 => x"2f",
  1437 => x"03",
  1438 => x"4e",
  1439 => x"95",
  1440 => x"2f",
  1441 => x"04",
  1442 => x"4e",
  1443 => x"95",
  1444 => x"20",
  1445 => x"0c",
  1446 => x"b1",
  1447 => x"87",
  1448 => x"84",
  1449 => x"87",
  1450 => x"4f",
  1451 => x"ef",
  1452 => x"00",
  1453 => x"10",
  1454 => x"2e",
  1455 => x"2a",
  1456 => x"00",
  1457 => x"08",
  1458 => x"bc",
  1459 => x"87",
  1460 => x"67",
  1461 => x"24",
  1462 => x"48",
  1463 => x"79",
  1464 => x"00",
  1465 => x"00",
  1466 => x"09",
  1467 => x"9c",
  1468 => x"4e",
  1469 => x"b9",
  1470 => x"00",
  1471 => x"00",
  1472 => x"08",
  1473 => x"06",
  1474 => x"2f",
  1475 => x"07",
  1476 => x"49",
  1477 => x"fa",
  1478 => x"fc",
  1479 => x"b2",
  1480 => x"4e",
  1481 => x"94",
  1482 => x"2f",
  1483 => x"03",
  1484 => x"4e",
  1485 => x"94",
  1486 => x"2f",
  1487 => x"04",
  1488 => x"4e",
  1489 => x"94",
  1490 => x"bd",
  1491 => x"87",
  1492 => x"84",
  1493 => x"87",
  1494 => x"4f",
  1495 => x"ef",
  1496 => x"00",
  1497 => x"10",
  1498 => x"2f",
  1499 => x"0b",
  1500 => x"4e",
  1501 => x"ba",
  1502 => x"fd",
  1503 => x"04",
  1504 => x"2e",
  1505 => x"2a",
  1506 => x"00",
  1507 => x"08",
  1508 => x"58",
  1509 => x"8f",
  1510 => x"bc",
  1511 => x"87",
  1512 => x"67",
  1513 => x"24",
  1514 => x"48",
  1515 => x"79",
  1516 => x"00",
  1517 => x"00",
  1518 => x"09",
  1519 => x"bf",
  1520 => x"4e",
  1521 => x"b9",
  1522 => x"00",
  1523 => x"00",
  1524 => x"08",
  1525 => x"06",
  1526 => x"2f",
  1527 => x"07",
  1528 => x"49",
  1529 => x"fa",
  1530 => x"fc",
  1531 => x"7e",
  1532 => x"4e",
  1533 => x"94",
  1534 => x"2f",
  1535 => x"03",
  1536 => x"4e",
  1537 => x"94",
  1538 => x"2f",
  1539 => x"04",
  1540 => x"4e",
  1541 => x"94",
  1542 => x"bf",
  1543 => x"86",
  1544 => x"84",
  1545 => x"86",
  1546 => x"4f",
  1547 => x"ef",
  1548 => x"00",
  1549 => x"10",
  1550 => x"2c",
  1551 => x"2a",
  1552 => x"00",
  1553 => x"0c",
  1554 => x"ba",
  1555 => x"86",
  1556 => x"67",
  1557 => x"24",
  1558 => x"48",
  1559 => x"79",
  1560 => x"00",
  1561 => x"00",
  1562 => x"09",
  1563 => x"e2",
  1564 => x"4e",
  1565 => x"b9",
  1566 => x"00",
  1567 => x"00",
  1568 => x"08",
  1569 => x"06",
  1570 => x"2f",
  1571 => x"06",
  1572 => x"49",
  1573 => x"fa",
  1574 => x"fc",
  1575 => x"52",
  1576 => x"4e",
  1577 => x"94",
  1578 => x"2f",
  1579 => x"03",
  1580 => x"4e",
  1581 => x"94",
  1582 => x"2f",
  1583 => x"04",
  1584 => x"4e",
  1585 => x"94",
  1586 => x"bb",
  1587 => x"86",
  1588 => x"84",
  1589 => x"86",
  1590 => x"4f",
  1591 => x"ef",
  1592 => x"00",
  1593 => x"10",
  1594 => x"2f",
  1595 => x"0b",
  1596 => x"4e",
  1597 => x"ba",
  1598 => x"fc",
  1599 => x"a4",
  1600 => x"2c",
  1601 => x"2a",
  1602 => x"00",
  1603 => x"0c",
  1604 => x"58",
  1605 => x"8f",
  1606 => x"ba",
  1607 => x"86",
  1608 => x"67",
  1609 => x"24",
  1610 => x"48",
  1611 => x"79",
  1612 => x"00",
  1613 => x"00",
  1614 => x"0a",
  1615 => x"05",
  1616 => x"4e",
  1617 => x"b9",
  1618 => x"00",
  1619 => x"00",
  1620 => x"08",
  1621 => x"06",
  1622 => x"2f",
  1623 => x"06",
  1624 => x"45",
  1625 => x"fa",
  1626 => x"fc",
  1627 => x"1e",
  1628 => x"4e",
  1629 => x"92",
  1630 => x"2f",
  1631 => x"03",
  1632 => x"4e",
  1633 => x"92",
  1634 => x"2f",
  1635 => x"04",
  1636 => x"4e",
  1637 => x"92",
  1638 => x"bd",
  1639 => x"85",
  1640 => x"84",
  1641 => x"85",
  1642 => x"4f",
  1643 => x"ef",
  1644 => x"00",
  1645 => x"10",
  1646 => x"20",
  1647 => x"02",
  1648 => x"4c",
  1649 => x"ee",
  1650 => x"3c",
  1651 => x"fc",
  1652 => x"ff",
  1653 => x"d8",
  1654 => x"4e",
  1655 => x"5e",
  1656 => x"4e",
  1657 => x"75",
  1658 => x"4e",
  1659 => x"56",
  1660 => x"00",
  1661 => x"00",
  1662 => x"48",
  1663 => x"e7",
  1664 => x"3f",
  1665 => x"30",
  1666 => x"2e",
  1667 => x"2e",
  1668 => x"00",
  1669 => x"08",
  1670 => x"48",
  1671 => x"79",
  1672 => x"00",
  1673 => x"00",
  1674 => x"0a",
  1675 => x"28",
  1676 => x"4e",
  1677 => x"b9",
  1678 => x"00",
  1679 => x"00",
  1680 => x"08",
  1681 => x"06",
  1682 => x"58",
  1683 => x"8f",
  1684 => x"42",
  1685 => x"83",
  1686 => x"42",
  1687 => x"82",
  1688 => x"47",
  1689 => x"fa",
  1690 => x"fd",
  1691 => x"0c",
  1692 => x"45",
  1693 => x"f9",
  1694 => x"00",
  1695 => x"00",
  1696 => x"07",
  1697 => x"e8",
  1698 => x"60",
  1699 => x"34",
  1700 => x"3f",
  1701 => x"04",
  1702 => x"42",
  1703 => x"67",
  1704 => x"2f",
  1705 => x"03",
  1706 => x"2f",
  1707 => x"07",
  1708 => x"4e",
  1709 => x"93",
  1710 => x"84",
  1711 => x"80",
  1712 => x"06",
  1713 => x"84",
  1714 => x"00",
  1715 => x"31",
  1716 => x"87",
  1717 => x"65",
  1718 => x"4f",
  1719 => x"ef",
  1720 => x"00",
  1721 => x"0c",
  1722 => x"0c",
  1723 => x"84",
  1724 => x"80",
  1725 => x"14",
  1726 => x"1f",
  1727 => x"2e",
  1728 => x"66",
  1729 => x"e2",
  1730 => x"48",
  1731 => x"78",
  1732 => x"00",
  1733 => x"2e",
  1734 => x"4e",
  1735 => x"92",
  1736 => x"06",
  1737 => x"83",
  1738 => x"00",
  1739 => x"21",
  1740 => x"23",
  1741 => x"45",
  1742 => x"58",
  1743 => x"8f",
  1744 => x"0c",
  1745 => x"83",
  1746 => x"80",
  1747 => x"05",
  1748 => x"41",
  1749 => x"91",
  1750 => x"67",
  1751 => x"04",
  1752 => x"42",
  1753 => x"84",
  1754 => x"60",
  1755 => x"c8",
  1756 => x"4a",
  1757 => x"82",
  1758 => x"67",
  1759 => x"18",
  1760 => x"48",
  1761 => x"79",
  1762 => x"00",
  1763 => x"00",
  1764 => x"0a",
  1765 => x"3d",
  1766 => x"4e",
  1767 => x"b9",
  1768 => x"00",
  1769 => x"00",
  1770 => x"08",
  1771 => x"06",
  1772 => x"2f",
  1773 => x"02",
  1774 => x"4e",
  1775 => x"ba",
  1776 => x"fb",
  1777 => x"88",
  1778 => x"50",
  1779 => x"8f",
  1780 => x"42",
  1781 => x"84",
  1782 => x"60",
  1783 => x"02",
  1784 => x"78",
  1785 => x"01",
  1786 => x"48",
  1787 => x"79",
  1788 => x"00",
  1789 => x"00",
  1790 => x"0a",
  1791 => x"5d",
  1792 => x"4e",
  1793 => x"b9",
  1794 => x"00",
  1795 => x"00",
  1796 => x"08",
  1797 => x"06",
  1798 => x"58",
  1799 => x"8f",
  1800 => x"42",
  1801 => x"85",
  1802 => x"42",
  1803 => x"83",
  1804 => x"47",
  1805 => x"fa",
  1806 => x"fc",
  1807 => x"18",
  1808 => x"45",
  1809 => x"f9",
  1810 => x"00",
  1811 => x"00",
  1812 => x"07",
  1813 => x"e8",
  1814 => x"60",
  1815 => x"32",
  1816 => x"2f",
  1817 => x"06",
  1818 => x"2f",
  1819 => x"05",
  1820 => x"2f",
  1821 => x"07",
  1822 => x"4e",
  1823 => x"93",
  1824 => x"86",
  1825 => x"80",
  1826 => x"06",
  1827 => x"86",
  1828 => x"00",
  1829 => x"19",
  1830 => x"87",
  1831 => x"65",
  1832 => x"4f",
  1833 => x"ef",
  1834 => x"00",
  1835 => x"0c",
  1836 => x"0c",
  1837 => x"86",
  1838 => x"80",
  1839 => x"0b",
  1840 => x"16",
  1841 => x"94",
  1842 => x"66",
  1843 => x"e4",
  1844 => x"48",
  1845 => x"78",
  1846 => x"00",
  1847 => x"2e",
  1848 => x"4e",
  1849 => x"92",
  1850 => x"06",
  1851 => x"85",
  1852 => x"00",
  1853 => x"13",
  1854 => x"45",
  1855 => x"67",
  1856 => x"58",
  1857 => x"8f",
  1858 => x"0c",
  1859 => x"85",
  1860 => x"80",
  1861 => x"0c",
  1862 => x"25",
  1863 => x"63",
  1864 => x"67",
  1865 => x"04",
  1866 => x"42",
  1867 => x"86",
  1868 => x"60",
  1869 => x"ca",
  1870 => x"4a",
  1871 => x"83",
  1872 => x"67",
  1873 => x"0a",
  1874 => x"2f",
  1875 => x"03",
  1876 => x"4e",
  1877 => x"ba",
  1878 => x"fb",
  1879 => x"22",
  1880 => x"58",
  1881 => x"8f",
  1882 => x"42",
  1883 => x"84",
  1884 => x"86",
  1885 => x"82",
  1886 => x"48",
  1887 => x"79",
  1888 => x"00",
  1889 => x"00",
  1890 => x"0a",
  1891 => x"77",
  1892 => x"4e",
  1893 => x"b9",
  1894 => x"00",
  1895 => x"00",
  1896 => x"08",
  1897 => x"06",
  1898 => x"58",
  1899 => x"8f",
  1900 => x"42",
  1901 => x"85",
  1902 => x"42",
  1903 => x"82",
  1904 => x"47",
  1905 => x"fa",
  1906 => x"fd",
  1907 => x"02",
  1908 => x"45",
  1909 => x"f9",
  1910 => x"00",
  1911 => x"00",
  1912 => x"07",
  1913 => x"e8",
  1914 => x"60",
  1915 => x"36",
  1916 => x"42",
  1917 => x"80",
  1918 => x"10",
  1919 => x"06",
  1920 => x"2f",
  1921 => x"00",
  1922 => x"2f",
  1923 => x"05",
  1924 => x"2f",
  1925 => x"07",
  1926 => x"4e",
  1927 => x"93",
  1928 => x"84",
  1929 => x"80",
  1930 => x"06",
  1931 => x"86",
  1932 => x"00",
  1933 => x"28",
  1934 => x"76",
  1935 => x"53",
  1936 => x"4f",
  1937 => x"ef",
  1938 => x"00",
  1939 => x"0c",
  1940 => x"0c",
  1941 => x"86",
  1942 => x"80",
  1943 => x"06",
  1944 => x"62",
  1945 => x"9e",
  1946 => x"66",
  1947 => x"e0",
  1948 => x"48",
  1949 => x"78",
  1950 => x"00",
  1951 => x"2e",
  1952 => x"4e",
  1953 => x"92",
  1954 => x"06",
  1955 => x"85",
  1956 => x"00",
  1957 => x"71",
  1958 => x"23",
  1959 => x"41",
  1960 => x"58",
  1961 => x"8f",
  1962 => x"0c",
  1963 => x"85",
  1964 => x"80",
  1965 => x"29",
  1966 => x"ef",
  1967 => x"a2",
  1968 => x"67",
  1969 => x"04",
  1970 => x"42",
  1971 => x"86",
  1972 => x"60",
  1973 => x"c6",
  1974 => x"4a",
  1975 => x"82",
  1976 => x"67",
  1977 => x"0a",
  1978 => x"2f",
  1979 => x"02",
  1980 => x"4e",
  1981 => x"ba",
  1982 => x"fa",
  1983 => x"ba",
  1984 => x"58",
  1985 => x"8f",
  1986 => x"42",
  1987 => x"84",
  1988 => x"84",
  1989 => x"83",
  1990 => x"67",
  1991 => x"14",
  1992 => x"48",
  1993 => x"79",
  1994 => x"00",
  1995 => x"00",
  1996 => x"0a",
  1997 => x"8c",
  1998 => x"4e",
  1999 => x"b9",
  2000 => x"00",
  2001 => x"00",
  2002 => x"08",
  2003 => x"06",
  2004 => x"2f",
  2005 => x"02",
  2006 => x"4e",
  2007 => x"ba",
  2008 => x"fa",
  2009 => x"a0",
  2010 => x"50",
  2011 => x"8f",
  2012 => x"20",
  2013 => x"04",
  2014 => x"4c",
  2015 => x"ee",
  2016 => x"0c",
  2017 => x"fc",
  2018 => x"ff",
  2019 => x"e0",
  2020 => x"4e",
  2021 => x"5e",
  2022 => x"4e",
  2023 => x"75",
  2024 => x"4e",
  2025 => x"56",
  2026 => x"00",
  2027 => x"00",
  2028 => x"20",
  2029 => x"2e",
  2030 => x"00",
  2031 => x"08",
  2032 => x"32",
  2033 => x"39",
  2034 => x"81",
  2035 => x"00",
  2036 => x"00",
  2037 => x"00",
  2038 => x"08",
  2039 => x"01",
  2040 => x"00",
  2041 => x"08",
  2042 => x"67",
  2043 => x"f4",
  2044 => x"33",
  2045 => x"c0",
  2046 => x"81",
  2047 => x"00",
  2048 => x"00",
  2049 => x"00",
  2050 => x"4e",
  2051 => x"5e",
  2052 => x"4e",
  2053 => x"75",
  2054 => x"4e",
  2055 => x"56",
  2056 => x"00",
  2057 => x"00",
  2058 => x"48",
  2059 => x"e7",
  2060 => x"20",
  2061 => x"30",
  2062 => x"24",
  2063 => x"6e",
  2064 => x"00",
  2065 => x"08",
  2066 => x"47",
  2067 => x"fa",
  2068 => x"ff",
  2069 => x"d4",
  2070 => x"60",
  2071 => x"0a",
  2072 => x"49",
  2073 => x"c0",
  2074 => x"2f",
  2075 => x"00",
  2076 => x"4e",
  2077 => x"93",
  2078 => x"52",
  2079 => x"82",
  2080 => x"58",
  2081 => x"8f",
  2082 => x"10",
  2083 => x"1a",
  2084 => x"66",
  2085 => x"f2",
  2086 => x"20",
  2087 => x"02",
  2088 => x"4c",
  2089 => x"ee",
  2090 => x"0c",
  2091 => x"04",
  2092 => x"ff",
  2093 => x"f4",
  2094 => x"4e",
  2095 => x"5e",
  2096 => x"4e",
  2097 => x"75",
  2098 => x"4d",
  2099 => x"69",
  2100 => x"73",
  2101 => x"61",
  2102 => x"6c",
  2103 => x"69",
  2104 => x"67",
  2105 => x"6e",
  2106 => x"65",
  2107 => x"64",
  2108 => x"20",
  2109 => x"6c",
  2110 => x"6f",
  2111 => x"6e",
  2112 => x"67",
  2113 => x"20",
  2114 => x"63",
  2115 => x"68",
  2116 => x"65",
  2117 => x"63",
  2118 => x"6b",
  2119 => x"20",
  2120 => x"28",
  2121 => x"63",
  2122 => x"61",
  2123 => x"63",
  2124 => x"68",
  2125 => x"65",
  2126 => x"29",
  2127 => x"20",
  2128 => x"66",
  2129 => x"61",
  2130 => x"69",
  2131 => x"6c",
  2132 => x"65",
  2133 => x"64",
  2134 => x"3a",
  2135 => x"20",
  2136 => x"00",
  2137 => x"4d",
  2138 => x"69",
  2139 => x"73",
  2140 => x"61",
  2141 => x"6c",
  2142 => x"69",
  2143 => x"67",
  2144 => x"6e",
  2145 => x"65",
  2146 => x"64",
  2147 => x"20",
  2148 => x"6c",
  2149 => x"6f",
  2150 => x"6e",
  2151 => x"67",
  2152 => x"20",
  2153 => x"63",
  2154 => x"68",
  2155 => x"65",
  2156 => x"63",
  2157 => x"6b",
  2158 => x"20",
  2159 => x"28",
  2160 => x"66",
  2161 => x"6c",
  2162 => x"75",
  2163 => x"73",
  2164 => x"68",
  2165 => x"29",
  2166 => x"20",
  2167 => x"66",
  2168 => x"61",
  2169 => x"69",
  2170 => x"6c",
  2171 => x"65",
  2172 => x"64",
  2173 => x"3a",
  2174 => x"20",
  2175 => x"00",
  2176 => x"4c",
  2177 => x"6f",
  2178 => x"6e",
  2179 => x"67",
  2180 => x"20",
  2181 => x"53",
  2182 => x"68",
  2183 => x"6f",
  2184 => x"72",
  2185 => x"74",
  2186 => x"20",
  2187 => x"63",
  2188 => x"68",
  2189 => x"65",
  2190 => x"63",
  2191 => x"6b",
  2192 => x"20",
  2193 => x"31",
  2194 => x"20",
  2195 => x"28",
  2196 => x"63",
  2197 => x"61",
  2198 => x"63",
  2199 => x"68",
  2200 => x"65",
  2201 => x"29",
  2202 => x"20",
  2203 => x"66",
  2204 => x"61",
  2205 => x"69",
  2206 => x"6c",
  2207 => x"65",
  2208 => x"64",
  2209 => x"3a",
  2210 => x"20",
  2211 => x"00",
  2212 => x"4c",
  2213 => x"6f",
  2214 => x"6e",
  2215 => x"67",
  2216 => x"20",
  2217 => x"53",
  2218 => x"68",
  2219 => x"6f",
  2220 => x"72",
  2221 => x"74",
  2222 => x"20",
  2223 => x"63",
  2224 => x"68",
  2225 => x"65",
  2226 => x"63",
  2227 => x"6b",
  2228 => x"20",
  2229 => x"31",
  2230 => x"20",
  2231 => x"28",
  2232 => x"66",
  2233 => x"6c",
  2234 => x"75",
  2235 => x"73",
  2236 => x"68",
  2237 => x"29",
  2238 => x"20",
  2239 => x"66",
  2240 => x"61",
  2241 => x"69",
  2242 => x"6c",
  2243 => x"65",
  2244 => x"64",
  2245 => x"3a",
  2246 => x"20",
  2247 => x"00",
  2248 => x"4c",
  2249 => x"6f",
  2250 => x"6e",
  2251 => x"67",
  2252 => x"20",
  2253 => x"53",
  2254 => x"68",
  2255 => x"6f",
  2256 => x"72",
  2257 => x"74",
  2258 => x"20",
  2259 => x"63",
  2260 => x"68",
  2261 => x"65",
  2262 => x"63",
  2263 => x"6b",
  2264 => x"20",
  2265 => x"32",
  2266 => x"20",
  2267 => x"28",
  2268 => x"63",
  2269 => x"61",
  2270 => x"63",
  2271 => x"68",
  2272 => x"65",
  2273 => x"29",
  2274 => x"20",
  2275 => x"66",
  2276 => x"61",
  2277 => x"69",
  2278 => x"6c",
  2279 => x"65",
  2280 => x"64",
  2281 => x"3a",
  2282 => x"20",
  2283 => x"00",
  2284 => x"4c",
  2285 => x"6f",
  2286 => x"6e",
  2287 => x"67",
  2288 => x"20",
  2289 => x"53",
  2290 => x"68",
  2291 => x"6f",
  2292 => x"72",
  2293 => x"74",
  2294 => x"20",
  2295 => x"63",
  2296 => x"68",
  2297 => x"65",
  2298 => x"63",
  2299 => x"6b",
  2300 => x"20",
  2301 => x"32",
  2302 => x"20",
  2303 => x"28",
  2304 => x"66",
  2305 => x"6c",
  2306 => x"75",
  2307 => x"73",
  2308 => x"68",
  2309 => x"29",
  2310 => x"20",
  2311 => x"66",
  2312 => x"61",
  2313 => x"69",
  2314 => x"6c",
  2315 => x"65",
  2316 => x"64",
  2317 => x"3a",
  2318 => x"20",
  2319 => x"00",
  2320 => x"4c",
  2321 => x"6f",
  2322 => x"6e",
  2323 => x"67",
  2324 => x"20",
  2325 => x"42",
  2326 => x"79",
  2327 => x"74",
  2328 => x"65",
  2329 => x"20",
  2330 => x"63",
  2331 => x"68",
  2332 => x"65",
  2333 => x"63",
  2334 => x"6b",
  2335 => x"20",
  2336 => x"31",
  2337 => x"20",
  2338 => x"28",
  2339 => x"63",
  2340 => x"61",
  2341 => x"63",
  2342 => x"68",
  2343 => x"65",
  2344 => x"29",
  2345 => x"20",
  2346 => x"66",
  2347 => x"61",
  2348 => x"69",
  2349 => x"6c",
  2350 => x"65",
  2351 => x"64",
  2352 => x"3a",
  2353 => x"20",
  2354 => x"00",
  2355 => x"4c",
  2356 => x"6f",
  2357 => x"6e",
  2358 => x"67",
  2359 => x"20",
  2360 => x"42",
  2361 => x"79",
  2362 => x"74",
  2363 => x"65",
  2364 => x"20",
  2365 => x"63",
  2366 => x"68",
  2367 => x"65",
  2368 => x"63",
  2369 => x"6b",
  2370 => x"20",
  2371 => x"31",
  2372 => x"20",
  2373 => x"28",
  2374 => x"66",
  2375 => x"6c",
  2376 => x"75",
  2377 => x"73",
  2378 => x"68",
  2379 => x"29",
  2380 => x"20",
  2381 => x"66",
  2382 => x"61",
  2383 => x"69",
  2384 => x"6c",
  2385 => x"65",
  2386 => x"64",
  2387 => x"3a",
  2388 => x"20",
  2389 => x"00",
  2390 => x"4c",
  2391 => x"6f",
  2392 => x"6e",
  2393 => x"67",
  2394 => x"20",
  2395 => x"42",
  2396 => x"79",
  2397 => x"74",
  2398 => x"65",
  2399 => x"20",
  2400 => x"63",
  2401 => x"68",
  2402 => x"65",
  2403 => x"63",
  2404 => x"6b",
  2405 => x"20",
  2406 => x"32",
  2407 => x"20",
  2408 => x"28",
  2409 => x"63",
  2410 => x"61",
  2411 => x"63",
  2412 => x"68",
  2413 => x"65",
  2414 => x"29",
  2415 => x"20",
  2416 => x"66",
  2417 => x"61",
  2418 => x"69",
  2419 => x"6c",
  2420 => x"65",
  2421 => x"64",
  2422 => x"3a",
  2423 => x"20",
  2424 => x"00",
  2425 => x"4c",
  2426 => x"6f",
  2427 => x"6e",
  2428 => x"67",
  2429 => x"20",
  2430 => x"42",
  2431 => x"79",
  2432 => x"74",
  2433 => x"65",
  2434 => x"20",
  2435 => x"63",
  2436 => x"68",
  2437 => x"65",
  2438 => x"63",
  2439 => x"6b",
  2440 => x"20",
  2441 => x"32",
  2442 => x"20",
  2443 => x"28",
  2444 => x"66",
  2445 => x"6c",
  2446 => x"75",
  2447 => x"73",
  2448 => x"68",
  2449 => x"29",
  2450 => x"20",
  2451 => x"66",
  2452 => x"61",
  2453 => x"69",
  2454 => x"6c",
  2455 => x"65",
  2456 => x"64",
  2457 => x"3a",
  2458 => x"20",
  2459 => x"00",
  2460 => x"4c",
  2461 => x"6f",
  2462 => x"6e",
  2463 => x"67",
  2464 => x"20",
  2465 => x"42",
  2466 => x"79",
  2467 => x"74",
  2468 => x"65",
  2469 => x"20",
  2470 => x"63",
  2471 => x"68",
  2472 => x"65",
  2473 => x"63",
  2474 => x"6b",
  2475 => x"20",
  2476 => x"33",
  2477 => x"20",
  2478 => x"28",
  2479 => x"63",
  2480 => x"61",
  2481 => x"63",
  2482 => x"68",
  2483 => x"65",
  2484 => x"29",
  2485 => x"20",
  2486 => x"66",
  2487 => x"61",
  2488 => x"69",
  2489 => x"6c",
  2490 => x"65",
  2491 => x"64",
  2492 => x"3a",
  2493 => x"20",
  2494 => x"00",
  2495 => x"4c",
  2496 => x"6f",
  2497 => x"6e",
  2498 => x"67",
  2499 => x"20",
  2500 => x"42",
  2501 => x"79",
  2502 => x"74",
  2503 => x"65",
  2504 => x"20",
  2505 => x"63",
  2506 => x"68",
  2507 => x"65",
  2508 => x"63",
  2509 => x"6b",
  2510 => x"20",
  2511 => x"33",
  2512 => x"20",
  2513 => x"28",
  2514 => x"66",
  2515 => x"6c",
  2516 => x"75",
  2517 => x"73",
  2518 => x"68",
  2519 => x"29",
  2520 => x"20",
  2521 => x"66",
  2522 => x"61",
  2523 => x"69",
  2524 => x"6c",
  2525 => x"65",
  2526 => x"64",
  2527 => x"3a",
  2528 => x"20",
  2529 => x"00",
  2530 => x"4c",
  2531 => x"6f",
  2532 => x"6e",
  2533 => x"67",
  2534 => x"20",
  2535 => x"42",
  2536 => x"79",
  2537 => x"74",
  2538 => x"65",
  2539 => x"20",
  2540 => x"63",
  2541 => x"68",
  2542 => x"65",
  2543 => x"63",
  2544 => x"6b",
  2545 => x"20",
  2546 => x"34",
  2547 => x"20",
  2548 => x"28",
  2549 => x"63",
  2550 => x"61",
  2551 => x"63",
  2552 => x"68",
  2553 => x"65",
  2554 => x"29",
  2555 => x"20",
  2556 => x"66",
  2557 => x"61",
  2558 => x"69",
  2559 => x"6c",
  2560 => x"65",
  2561 => x"64",
  2562 => x"3a",
  2563 => x"20",
  2564 => x"00",
  2565 => x"4c",
  2566 => x"6f",
  2567 => x"6e",
  2568 => x"67",
  2569 => x"20",
  2570 => x"42",
  2571 => x"79",
  2572 => x"74",
  2573 => x"65",
  2574 => x"20",
  2575 => x"63",
  2576 => x"68",
  2577 => x"65",
  2578 => x"63",
  2579 => x"6b",
  2580 => x"20",
  2581 => x"34",
  2582 => x"20",
  2583 => x"28",
  2584 => x"66",
  2585 => x"6c",
  2586 => x"75",
  2587 => x"73",
  2588 => x"68",
  2589 => x"29",
  2590 => x"20",
  2591 => x"66",
  2592 => x"61",
  2593 => x"69",
  2594 => x"6c",
  2595 => x"65",
  2596 => x"64",
  2597 => x"3a",
  2598 => x"20",
  2599 => x"00",
  2600 => x"0a",
  2601 => x"4c",
  2602 => x"6f",
  2603 => x"6e",
  2604 => x"67",
  2605 => x"2f",
  2606 => x"73",
  2607 => x"68",
  2608 => x"6f",
  2609 => x"72",
  2610 => x"74",
  2611 => x"20",
  2612 => x"74",
  2613 => x"65",
  2614 => x"73",
  2615 => x"74",
  2616 => x"2e",
  2617 => x"2e",
  2618 => x"2e",
  2619 => x"0a",
  2620 => x"00",
  2621 => x"42",
  2622 => x"61",
  2623 => x"64",
  2624 => x"20",
  2625 => x"62",
  2626 => x"69",
  2627 => x"74",
  2628 => x"73",
  2629 => x"20",
  2630 => x"66",
  2631 => x"72",
  2632 => x"6f",
  2633 => x"6d",
  2634 => x"20",
  2635 => x"4c",
  2636 => x"6f",
  2637 => x"6e",
  2638 => x"67",
  2639 => x"20",
  2640 => x"53",
  2641 => x"68",
  2642 => x"6f",
  2643 => x"72",
  2644 => x"74",
  2645 => x"20",
  2646 => x"74",
  2647 => x"65",
  2648 => x"73",
  2649 => x"74",
  2650 => x"3a",
  2651 => x"20",
  2652 => x"00",
  2653 => x"0a",
  2654 => x"4d",
  2655 => x"69",
  2656 => x"73",
  2657 => x"61",
  2658 => x"6c",
  2659 => x"69",
  2660 => x"67",
  2661 => x"6e",
  2662 => x"65",
  2663 => x"64",
  2664 => x"20",
  2665 => x"4c",
  2666 => x"6f",
  2667 => x"6e",
  2668 => x"67",
  2669 => x"20",
  2670 => x"74",
  2671 => x"65",
  2672 => x"73",
  2673 => x"74",
  2674 => x"2e",
  2675 => x"2e",
  2676 => x"2e",
  2677 => x"0a",
  2678 => x"00",
  2679 => x"4c",
  2680 => x"6f",
  2681 => x"6e",
  2682 => x"67",
  2683 => x"20",
  2684 => x"2f",
  2685 => x"20",
  2686 => x"62",
  2687 => x"79",
  2688 => x"74",
  2689 => x"65",
  2690 => x"20",
  2691 => x"74",
  2692 => x"65",
  2693 => x"73",
  2694 => x"74",
  2695 => x"2e",
  2696 => x"2e",
  2697 => x"2e",
  2698 => x"0a",
  2699 => x"00",
  2700 => x"42",
  2701 => x"61",
  2702 => x"64",
  2703 => x"20",
  2704 => x"62",
  2705 => x"69",
  2706 => x"74",
  2707 => x"73",
  2708 => x"20",
  2709 => x"64",
  2710 => x"65",
  2711 => x"74",
  2712 => x"65",
  2713 => x"63",
  2714 => x"74",
  2715 => x"65",
  2716 => x"64",
  2717 => x"3a",
  2718 => x"20",
  2719 => x"00",
  2720 => x"43",
  2721 => x"6f",
  2722 => x"6d",
  2723 => x"6d",
  2724 => x"65",
  2725 => x"6e",
  2726 => x"63",
  2727 => x"69",
  2728 => x"6e",
  2729 => x"67",
  2730 => x"20",
  2731 => x"73",
  2732 => x"61",
  2733 => x"6e",
  2734 => x"69",
  2735 => x"74",
  2736 => x"79",
  2737 => x"20",
  2738 => x"63",
  2739 => x"68",
  2740 => x"65",
  2741 => x"63",
  2742 => x"6b",
  2743 => x"73",
  2744 => x"2e",
  2745 => x"2e",
  2746 => x"2e",
  2747 => x"0a",
  2748 => x"00",
  2749 => x"4d",
  2750 => x"65",
  2751 => x"6d",
  2752 => x"6f",
  2753 => x"72",
  2754 => x"79",
  2755 => x"20",
  2756 => x"63",
  2757 => x"68",
  2758 => x"65",
  2759 => x"63",
  2760 => x"6b",
  2761 => x"20",
  2762 => x"70",
  2763 => x"61",
  2764 => x"73",
  2765 => x"73",
  2766 => x"65",
  2767 => x"64",
  2768 => x"0a",
  2769 => x"00",
  2770 => x"4d",
  2771 => x"65",
  2772 => x"6d",
  2773 => x"6f",
  2774 => x"72",
  2775 => x"79",
  2776 => x"20",
  2777 => x"63",
  2778 => x"68",
  2779 => x"65",
  2780 => x"63",
  2781 => x"6b",
  2782 => x"20",
  2783 => x"66",
  2784 => x"61",
  2785 => x"69",
  2786 => x"6c",
  2787 => x"65",
  2788 => x"64",
  2789 => x"0a",
  2790 => x"00",
  2791 => x"00",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;

