
--
-- Copyright (c) 2008-2019 Sytse van Slooten
--
-- Permission is hereby granted to any person obtaining a copy of these VHDL source files and
-- other language source files and associated documentation files ("the materials") to use
-- these materials solely for personal, non-commercial purposes.
-- You are also granted permission to make changes to the materials, on the condition that this
-- copyright notice is retained unchanged.
--
-- The materials are distributed in the hope that they will be useful, but WITHOUT ANY WARRANTY;
-- without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
--

-- $Revision: 1.8 $

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity blockram2 is
   port(
      base_addr : in std_logic_vector(17 downto 0);

      bus_addr_match : out std_logic;
      bus_addr : in std_logic_vector(17 downto 0);
      bus_dati : out std_logic_vector(15 downto 0);
      bus_dato : in std_logic_vector(15 downto 0);
      bus_control_dati : in std_logic;
      bus_control_dato : in std_logic;
      bus_control_datob : in std_logic;

      reset : in std_logic;
      clk : in std_logic
   );
end blockram2;

architecture implementation of blockram2 is

signal base_addr_match : std_logic;

subtype u is std_logic_vector(7 downto 0);
type mem_type is array(0 to 2047) of u;

-- code base at 130000

signal meme : mem_type := mem_type'(
u'(x"5f"),u'(x"72"),u'(x"4f"),u'(x"54"),u'(x"31"),u'(x"df"),u'(x"d2"),u'(x"0c"),u'(x"df"),u'(x"e0"),u'(x"0e"),u'(x"c6"),u'(x"8a"),u'(x"80"),u'(x"01"),u'(x"26"),
u'(x"d0"),u'(x"ff"),u'(x"97"),u'(x"6a"),u'(x"fa"),u'(x"df"),u'(x"00"),u'(x"76"),u'(x"1f"),u'(x"dc"),u'(x"1f"),u'(x"da"),u'(x"df"),u'(x"07"),u'(x"7c"),u'(x"5f"),
u'(x"3c"),u'(x"00"),u'(x"80"),u'(x"c4"),u'(x"40"),u'(x"fc"),u'(x"c4"),u'(x"40"),u'(x"e6"),u'(x"20"),u'(x"c0"),u'(x"08"),u'(x"ce"),u'(x"c0"),u'(x"1b"),u'(x"04"),
u'(x"ce"),u'(x"24"),u'(x"c0"),u'(x"f8"),u'(x"80"),u'(x"5f"),u'(x"1a"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"c4"),u'(x"00"),u'(x"c4"),u'(x"c4"),u'(x"04"),u'(x"82"),
u'(x"87"),u'(x"5f"),u'(x"48"),u'(x"c1"),u'(x"20"),u'(x"01"),u'(x"13"),u'(x"4c"),u'(x"17"),u'(x"41"),u'(x"0b"),u'(x"c1"),u'(x"09"),u'(x"17"),u'(x"24"),u'(x"0a"),
u'(x"17"),u'(x"2e"),u'(x"41"),u'(x"17"),u'(x"39"),u'(x"02"),u'(x"17"),u'(x"5a"),u'(x"3b"),u'(x"40"),u'(x"40"),u'(x"dc"),u'(x"11"),u'(x"07"),u'(x"c9"),u'(x"fc"),
u'(x"c0"),u'(x"38"),u'(x"c0"),u'(x"08"),u'(x"67"),u'(x"87"),u'(x"c0"),u'(x"d4"),u'(x"df"),u'(x"d8"),u'(x"14"),u'(x"c0"),u'(x"8a"),u'(x"c3"),u'(x"03"),u'(x"c5"),
u'(x"c2"),u'(x"06"),u'(x"c2"),u'(x"70"),u'(x"c4"),u'(x"74"),u'(x"8a"),u'(x"6f"),u'(x"50"),u'(x"17"),u'(x"9a"),u'(x"fc"),u'(x"6a"),u'(x"c0"),u'(x"d4"),u'(x"d7"),
u'(x"d2"),u'(x"02"),u'(x"49"),u'(x"66"),u'(x"c5"),u'(x"d8"),u'(x"c4"),u'(x"c4"),u'(x"8a"),u'(x"26"),u'(x"5f"),u'(x"36"),u'(x"c2"),u'(x"02"),u'(x"5f"),u'(x"96"),
u'(x"3b"),u'(x"00"),u'(x"5f"),u'(x"b0"),u'(x"d6"),u'(x"64"),u'(x"5f"),u'(x"8a"),u'(x"5f"),u'(x"36"),u'(x"84"),u'(x"c3"),u'(x"04"),u'(x"df"),u'(x"42"),u'(x"c3"),
u'(x"fc"),u'(x"02"),u'(x"df"),u'(x"82"),u'(x"97"),u'(x"03"),u'(x"fb"),u'(x"5f"),u'(x"a6"),u'(x"20"),u'(x"4b"),u'(x"5f"),u'(x"48"),u'(x"c1"),u'(x"f0"),u'(x"df"),
u'(x"b8"),u'(x"04"),u'(x"03"),u'(x"c1"),u'(x"e9"),u'(x"44"),u'(x"82"),u'(x"c4"),u'(x"c4"),u'(x"6a"),u'(x"17"),u'(x"8a"),u'(x"02"),u'(x"c4"),u'(x"9a"),u'(x"5f"),
u'(x"a6"),u'(x"2f"),u'(x"73"),u'(x"df"),u'(x"dc"),u'(x"df"),u'(x"02"),u'(x"d2"),u'(x"03"),u'(x"c2"),u'(x"d4"),u'(x"85"),u'(x"17"),u'(x"9f"),u'(x"da"),u'(x"17"),
u'(x"5f"),u'(x"86"),u'(x"82"),u'(x"0a"),u'(x"5f"),u'(x"86"),u'(x"81"),u'(x"81"),u'(x"c1"),u'(x"42"),u'(x"03"),u'(x"5f"),u'(x"86"),u'(x"82"),u'(x"df"),u'(x"d4"),
u'(x"d6"),u'(x"9f"),u'(x"d4"),u'(x"7f"),u'(x"5f"),u'(x"a6"),u'(x"3f"),u'(x"1f"),u'(x"d2"),u'(x"5f"),u'(x"a2"),u'(x"2a"),u'(x"1f"),u'(x"d8"),u'(x"03"),u'(x"05"),
u'(x"1f"),u'(x"d0"),u'(x"1f"),u'(x"dd"),u'(x"04"),u'(x"02"),u'(x"c6"),u'(x"6a"),u'(x"5f"),u'(x"48"),u'(x"17"),u'(x"2d"),u'(x"05"),u'(x"c2"),u'(x"e5"),u'(x"9f"),
u'(x"dd"),u'(x"f4"),u'(x"c1"),u'(x"fb"),u'(x"df"),u'(x"b8"),u'(x"04"),u'(x"c4"),u'(x"df"),u'(x"78"),u'(x"eb"),u'(x"9f"),u'(x"dd"),u'(x"01"),u'(x"04"),u'(x"c4"),
u'(x"d0"),u'(x"c1"),u'(x"79"),u'(x"c2"),u'(x"c2"),u'(x"ce"),u'(x"c4"),u'(x"d0"),u'(x"c4"),u'(x"02"),u'(x"8a"),u'(x"9f"),u'(x"d0"),u'(x"82"),u'(x"d1"),u'(x"d2"),
u'(x"83"),u'(x"05"),u'(x"9f"),u'(x"d8"),u'(x"cb"),u'(x"c3"),u'(x"0b"),u'(x"5f"),u'(x"84"),u'(x"5f"),u'(x"36"),u'(x"df"),u'(x"02"),u'(x"d2"),u'(x"40"),u'(x"5f"),
u'(x"c4"),u'(x"b5"),u'(x"c4"),u'(x"84"),u'(x"c2"),u'(x"c0"),u'(x"df"),u'(x"02"),u'(x"d2"),u'(x"04"),u'(x"44"),u'(x"df"),u'(x"01"),u'(x"d2"),u'(x"c2"),u'(x"02"),
u'(x"1f"),u'(x"d4"),u'(x"c4"),u'(x"d4"),u'(x"df"),u'(x"01"),u'(x"d2"),u'(x"05"),u'(x"84"),u'(x"f0"),u'(x"c0"),u'(x"d4"),u'(x"01"),u'(x"00"),u'(x"5f"),u'(x"c4"),
u'(x"9b"),u'(x"df"),u'(x"dc"),u'(x"93"),u'(x"9f"),u'(x"d9"),u'(x"c0"),u'(x"d2"),u'(x"8b"),u'(x"df"),u'(x"dc"),u'(x"df"),u'(x"d9"),u'(x"03"),u'(x"df"),u'(x"d6"),
u'(x"d4"),u'(x"1f"),u'(x"d4"),u'(x"5f"),u'(x"26"),u'(x"e6"),u'(x"d2"),u'(x"df"),u'(x"02"),u'(x"d2"),u'(x"c0"),u'(x"d4"),u'(x"5f"),u'(x"8e"),u'(x"9f"),u'(x"d2"),
u'(x"c0"),u'(x"5c"),u'(x"d6"),u'(x"01"),u'(x"c0"),u'(x"5f"),u'(x"1a"),u'(x"ca"),u'(x"c0"),u'(x"d2"),u'(x"dd"),u'(x"df"),u'(x"dc"),u'(x"1f"),u'(x"d4"),u'(x"e3"),
u'(x"c0"),u'(x"18"),u'(x"c4"),u'(x"c3"),u'(x"11"),u'(x"85"),u'(x"7a"),u'(x"c5"),u'(x"c4"),u'(x"9a"),u'(x"c2"),u'(x"08"),u'(x"74"),u'(x"0c"),u'(x"05"),u'(x"17"),
u'(x"a8"),u'(x"6f"),u'(x"d4"),u'(x"f9"),u'(x"4c"),u'(x"bd"),u'(x"c2"),u'(x"06"),u'(x"68"),u'(x"34"),u'(x"9a"),u'(x"34"),u'(x"ac"),u'(x"b5"),u'(x"04"),u'(x"f4"),
u'(x"18"),u'(x"9a"),u'(x"f4"),u'(x"d2"),u'(x"be"),u'(x"34"),u'(x"ac"),u'(x"d4"),u'(x"17"),u'(x"10"),u'(x"f4"),u'(x"a7"),u'(x"df"),u'(x"02"),u'(x"d2"),u'(x"51"),
u'(x"5f"),u'(x"a6"),u'(x"20"),u'(x"c3"),u'(x"4c"),u'(x"c5"),u'(x"d4"),u'(x"c5"),u'(x"c5"),u'(x"40"),u'(x"5f"),u'(x"c4"),u'(x"40"),u'(x"80"),u'(x"0c"),u'(x"c0"),
u'(x"80"),u'(x"09"),u'(x"c0"),u'(x"7f"),u'(x"06"),u'(x"df"),u'(x"d2"),u'(x"5f"),u'(x"c4"),u'(x"9f"),u'(x"d2"),u'(x"5f"),u'(x"d8"),u'(x"c0"),u'(x"80"),u'(x"01"),
u'(x"02"),u'(x"00"),u'(x"42"),u'(x"d7"),u'(x"4d"),u'(x"81"),u'(x"01"),u'(x"01"),u'(x"c3"),u'(x"27"),u'(x"df"),u'(x"02"),u'(x"d2"),u'(x"c2"),u'(x"80"),u'(x"c4"),
u'(x"7e"),u'(x"44"),u'(x"9f"),u'(x"82"),u'(x"c6"),u'(x"df"),u'(x"70"),u'(x"c3"),u'(x"e6"),u'(x"2f"),u'(x"80"),u'(x"c1"),u'(x"1e"),u'(x"00"),u'(x"05"),u'(x"05"),
u'(x"0e"),u'(x"26"),u'(x"5f"),u'(x"26"),u'(x"80"),u'(x"5f"),u'(x"8e"),u'(x"80"),u'(x"02"),u'(x"5f"),u'(x"1a"),u'(x"80"),u'(x"5f"),u'(x"c4"),u'(x"84"),u'(x"96"),
u'(x"e1"),u'(x"5f"),u'(x"c8"),u'(x"5f"),u'(x"9a"),u'(x"11"),u'(x"cb"),u'(x"5f"),u'(x"9a"),u'(x"11"),u'(x"c7"),u'(x"ce"),u'(x"05"),u'(x"e2"),u'(x"ce"),u'(x"5f"),
u'(x"03"),u'(x"83"),u'(x"83"),u'(x"83"),u'(x"c5"),u'(x"da"),u'(x"ce"),u'(x"00"),u'(x"80"),u'(x"c0"),u'(x"80"),u'(x"05"),u'(x"d3"),u'(x"c3"),u'(x"e2"),u'(x"df"),
u'(x"11"),u'(x"dc"),u'(x"85"),u'(x"dd"),u'(x"c5"),u'(x"5f"),u'(x"78"),u'(x"5f"),u'(x"b0"),u'(x"1f"),u'(x"db"),u'(x"df"),u'(x"da"),u'(x"0b"),u'(x"c4"),u'(x"0e"),
u'(x"34"),u'(x"9a"),u'(x"be"),u'(x"fc"),u'(x"03"),u'(x"9a"),u'(x"c4"),u'(x"c4"),u'(x"f7"),u'(x"80"),u'(x"81"),u'(x"82"),u'(x"83"),u'(x"84"),u'(x"85"),u'(x"86"),
u'(x"e6"),u'(x"7a"),u'(x"ce"),u'(x"10"),u'(x"9f"),u'(x"fe"),u'(x"df"),u'(x"da"),u'(x"08"),u'(x"ce"),u'(x"10"),u'(x"df"),u'(x"d2"),u'(x"0c"),u'(x"df"),u'(x"e0"),
u'(x"0e"),u'(x"e6"),u'(x"78"),u'(x"06"),u'(x"c0"),u'(x"dc"),u'(x"aa"),u'(x"c2"),u'(x"a8"),u'(x"c3"),u'(x"02"),u'(x"70"),u'(x"ac"),u'(x"5f"),u'(x"b0"),u'(x"d7"),
u'(x"dc"),u'(x"0e"),u'(x"c6"),u'(x"df"),u'(x"da"),u'(x"c3"),u'(x"9f"),u'(x"db"),u'(x"d0"),u'(x"9f"),u'(x"78"),u'(x"9f"),u'(x"7a"),u'(x"df"),u'(x"11"),u'(x"dc"),
u'(x"9f"),u'(x"76"),u'(x"c6"),u'(x"76"),u'(x"66"),u'(x"26"),u'(x"e6"),u'(x"a6"),u'(x"66"),u'(x"26"),u'(x"c4"),u'(x"db"),u'(x"05"),u'(x"c4"),u'(x"aa"),u'(x"5f"),
u'(x"a2"),u'(x"23"),u'(x"df"),u'(x"da"),u'(x"08"),u'(x"04"),u'(x"3c"),u'(x"be"),u'(x"9a"),u'(x"d4"),u'(x"17"),u'(x"0e"),u'(x"f9"),u'(x"c5"),u'(x"78"),u'(x"df"),
u'(x"da"),u'(x"14"),u'(x"e5"),u'(x"5f"),u'(x"78"),u'(x"c4"),u'(x"0e"),u'(x"74"),u'(x"9a"),u'(x"10"),u'(x"c4"),u'(x"c4"),u'(x"fa"),u'(x"5f"),u'(x"72"),u'(x"42"),
u'(x"20"),u'(x"40"),u'(x"df"),u'(x"02"),u'(x"78"),u'(x"1a"),u'(x"c4"),u'(x"10"),u'(x"74"),u'(x"9a"),u'(x"1f"),u'(x"dc"),u'(x"f4"),u'(x"ac"),u'(x"b0"),u'(x"f4"),
u'(x"01"),u'(x"ac"),u'(x"5f"),u'(x"72"),u'(x"42"),u'(x"c0"),u'(x"dc"),u'(x"80"),u'(x"c0"),u'(x"30"),u'(x"5f"),u'(x"30"),u'(x"c4"),u'(x"dc"),u'(x"00"),u'(x"9a"),
u'(x"df"),u'(x"02"),u'(x"d2"),u'(x"5f"),u'(x"8e"),u'(x"5f"),u'(x"ce"),u'(x"df"),u'(x"88"),u'(x"18"),u'(x"26"),u'(x"c4"),u'(x"8a"),u'(x"c0"),u'(x"16"),u'(x"8c"),
u'(x"03"),u'(x"08"),u'(x"01"),u'(x"00"),u'(x"d4"),u'(x"17"),u'(x"9a"),u'(x"f7"),u'(x"0e"),u'(x"c0"),u'(x"8a"),u'(x"05"),u'(x"80"),u'(x"c0"),u'(x"30"),u'(x"5f"),
u'(x"30"),u'(x"80"),u'(x"c3"),u'(x"06"),u'(x"c4"),u'(x"fe"),u'(x"df"),u'(x"01"),u'(x"d2"),u'(x"13"),u'(x"26"),u'(x"83"),u'(x"84"),u'(x"c0"),u'(x"5f"),u'(x"fa"),
u'(x"5f"),u'(x"36"),u'(x"ce"),u'(x"80"),u'(x"97"),u'(x"20"),u'(x"02"),u'(x"ce"),u'(x"3f"),u'(x"c0"),u'(x"00"),u'(x"80"),u'(x"1b"),u'(x"26"),u'(x"c4"),u'(x"03"),
u'(x"00"),u'(x"4e"),u'(x"40"),u'(x"c4"),u'(x"fc"),u'(x"c0"),u'(x"30"),u'(x"5f"),u'(x"1a"),u'(x"c3"),u'(x"f3"),u'(x"d6"),u'(x"c0"),u'(x"df"),u'(x"74"),u'(x"fd"),
u'(x"1f"),u'(x"76"),u'(x"85"),u'(x"c0"),u'(x"0d"),u'(x"5f"),u'(x"30"),u'(x"00"),u'(x"5f"),u'(x"1a"),u'(x"f1"),u'(x"c0"),u'(x"3d"),u'(x"ef"),u'(x"df"),u'(x"70"),
u'(x"fd"),u'(x"c0"),u'(x"72"),u'(x"87"),u'(x"df"),u'(x"3c"),u'(x"80"),u'(x"c0"),u'(x"80"),u'(x"c0"),u'(x"f9"),u'(x"17"),u'(x"0a"),u'(x"0a"),u'(x"17"),u'(x"60"),
u'(x"02"),u'(x"c0"),u'(x"20"),u'(x"5f"),u'(x"1a"),u'(x"c0"),u'(x"20"),u'(x"ec"),u'(x"85"),u'(x"c0"),u'(x"7c"),u'(x"03"),u'(x"c0"),u'(x"7a"),u'(x"04"),u'(x"80"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"c0"),u'(x"10"),u'(x"1f"),u'(x"fe"),u'(x"df"),u'(x"70"),u'(x"de"),u'(x"df"),u'(x"74"),u'(x"df"),u'(x"1f"),u'(x"70"),u'(x"1f"),
u'(x"74"),u'(x"5f"),u'(x"26"),u'(x"40"),u'(x"bd"),u'(x"5f"),u'(x"1a"),u'(x"fb"),u'(x"df"),u'(x"e0"),u'(x"fe"),u'(x"5f"),u'(x"26"),u'(x"df"),u'(x"74"),u'(x"fd"),
u'(x"df"),u'(x"00"),u'(x"70"),u'(x"03"),u'(x"df"),u'(x"70"),u'(x"fd"),u'(x"df"),u'(x"de"),u'(x"70"),u'(x"df"),u'(x"df"),u'(x"74"),u'(x"85"),u'(x"c2"),u'(x"0a"),
u'(x"df"),u'(x"01"),u'(x"d2"),u'(x"04"),u'(x"05"),u'(x"3f"),u'(x"d4"),u'(x"02"),u'(x"3f"),u'(x"d4"),u'(x"87"),u'(x"df"),u'(x"3c"),u'(x"e6"),u'(x"04"),u'(x"4e"),
u'(x"02"),u'(x"ce"),u'(x"86"),u'(x"c5"),u'(x"3c"),u'(x"01"),u'(x"03"),u'(x"cd"),u'(x"c0"),u'(x"fc"),u'(x"cd"),u'(x"df"),u'(x"50"),u'(x"02"),u'(x"c2"),u'(x"04"),
u'(x"df"),u'(x"50"),u'(x"84"),u'(x"c2"),u'(x"19"),u'(x"01"),u'(x"cd"),u'(x"04"),u'(x"c3"),u'(x"ec"),u'(x"03"),u'(x"ea"),u'(x"11"),u'(x"f8"),u'(x"df"),u'(x"01"),
u'(x"70"),u'(x"df"),u'(x"3c"),u'(x"c0"),u'(x"00"),u'(x"03"),u'(x"c2"),u'(x"87"),u'(x"cd"),u'(x"04"),u'(x"cd"),u'(x"c0"),u'(x"04"),u'(x"87"),u'(x"82"),u'(x"81"),
u'(x"81"),u'(x"5f"),u'(x"86"),u'(x"cd"),u'(x"c3"),u'(x"e4"),u'(x"84"),u'(x"1f"),u'(x"78"),u'(x"df"),u'(x"11"),u'(x"dc"),u'(x"5f"),u'(x"ce"),u'(x"df"),u'(x"3c"),
u'(x"c3"),u'(x"ae"),u'(x"01"),u'(x"00"),u'(x"80"),u'(x"4b"),u'(x"00"),u'(x"c0"),u'(x"06"),u'(x"40"),u'(x"4b"),u'(x"40"),u'(x"4b"),u'(x"44"),u'(x"04"),u'(x"40"),
u'(x"5f"),u'(x"b4"),u'(x"fa"),u'(x"40"),u'(x"4b"),u'(x"4b"),u'(x"e5"),u'(x"5f"),u'(x"b4"),u'(x"c0"),u'(x"01"),u'(x"5f"),u'(x"1a"),u'(x"ac"),u'(x"a2"),u'(x"fa"),
u'(x"56"),u'(x"28"),u'(x"6c"),u'(x"40"),u'(x"a8"),u'(x"a8"),u'(x"a0"),u'(x"00"),u'(x"4a"),u'(x"7c"),u'(x"aa"),u'(x"0e"),u'(x"3a"),u'(x"06"),u'(x"f6"),u'(x"58"),
u'(x"a8"),u'(x"cc"),u'(x"9a"),u'(x"ae"),u'(x"2c"),u'(x"76"),u'(x"f0"),u'(x"b6"),u'(x"53"),u'(x"4d"),u'(x"55"),u'(x"41"),u'(x"52"),u'(x"00"),u'(x"0d"),u'(x"24"),
u'(x"2f"),u'(x"3c"),u'(x"40"),u'(x"43"),u'(x"45"),u'(x"47"),u'(x"4c"),u'(x"50"),u'(x"53"),u'(x"58"),u'(x"5e"),u'(x"00"),u'(x"03"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00") 
);
signal memo : mem_type := mem_type'(
u'(x"09"),u'(x"b6"),u'(x"44"),u'(x"31"),u'(x"00"),u'(x"15"),u'(x"b4"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"b8"),u'(x"11"),u'(x"0a"),u'(x"0a"),
u'(x"15"),u'(x"ff"),u'(x"21"),u'(x"b8"),u'(x"82"),u'(x"15"),u'(x"02"),u'(x"b8"),u'(x"98"),u'(x"b8"),u'(x"0a"),u'(x"b8"),u'(x"15"),u'(x"00"),u'(x"b8"),u'(x"00"),
u'(x"b3"),u'(x"0a"),u'(x"0a"),u'(x"e5"),u'(x"06"),u'(x"86"),u'(x"65"),u'(x"06"),u'(x"15"),u'(x"5b"),u'(x"0a"),u'(x"03"),u'(x"00"),u'(x"e5"),u'(x"00"),u'(x"87"),
u'(x"15"),u'(x"48"),u'(x"0b"),u'(x"02"),u'(x"65"),u'(x"09"),u'(x"b6"),u'(x"0a"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"61"),u'(x"0c"),u'(x"0c"),u'(x"60"),u'(x"0a"),
u'(x"00"),u'(x"09"),u'(x"b6"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"03"),u'(x"87"),u'(x"20"),u'(x"00"),u'(x"86"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"00"),u'(x"03"),
u'(x"20"),u'(x"00"),u'(x"87"),u'(x"20"),u'(x"00"),u'(x"01"),u'(x"20"),u'(x"00"),u'(x"82"),u'(x"e0"),u'(x"e0"),u'(x"01"),u'(x"a0"),u'(x"03"),u'(x"8b"),u'(x"02"),
u'(x"e5"),u'(x"00"),u'(x"65"),u'(x"00"),u'(x"86"),u'(x"00"),u'(x"17"),u'(x"b8"),u'(x"8b"),u'(x"b8"),u'(x"03"),u'(x"15"),u'(x"b8"),u'(x"0a"),u'(x"80"),u'(x"10"),
u'(x"0b"),u'(x"03"),u'(x"0a"),u'(x"06"),u'(x"0c"),u'(x"11"),u'(x"b8"),u'(x"01"),u'(x"11"),u'(x"20"),u'(x"b8"),u'(x"87"),u'(x"01"),u'(x"15"),u'(x"b8"),u'(x"27"),
u'(x"b8"),u'(x"00"),u'(x"02"),u'(x"11"),u'(x"15"),u'(x"b1"),u'(x"0c"),u'(x"65"),u'(x"b8"),u'(x"12"),u'(x"09"),u'(x"b6"),u'(x"0a"),u'(x"80"),u'(x"00"),u'(x"b5"),
u'(x"02"),u'(x"11"),u'(x"00"),u'(x"b5"),u'(x"0b"),u'(x"01"),u'(x"09"),u'(x"b1"),u'(x"09"),u'(x"b6"),u'(x"12"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"b0"),u'(x"0a"),
u'(x"02"),u'(x"0a"),u'(x"09"),u'(x"b0"),u'(x"20"),u'(x"00"),u'(x"87"),u'(x"09"),u'(x"b6"),u'(x"00"),u'(x"01"),u'(x"09"),u'(x"b6"),u'(x"15"),u'(x"b7"),u'(x"09"),
u'(x"b0"),u'(x"10"),u'(x"87"),u'(x"e5"),u'(x"b7"),u'(x"10"),u'(x"0a"),u'(x"0c"),u'(x"65"),u'(x"b8"),u'(x"21"),u'(x"b8"),u'(x"83"),u'(x"15"),u'(x"b8"),u'(x"09"),
u'(x"b6"),u'(x"00"),u'(x"01"),u'(x"09"),u'(x"b6"),u'(x"25"),u'(x"00"),u'(x"b8"),u'(x"02"),u'(x"17"),u'(x"b8"),u'(x"00"),u'(x"01"),u'(x"90"),u'(x"b8"),u'(x"01"),
u'(x"09"),u'(x"b1"),u'(x"12"),u'(x"01"),u'(x"09"),u'(x"b1"),u'(x"92"),u'(x"0a"),u'(x"0c"),u'(x"60"),u'(x"01"),u'(x"09"),u'(x"b1"),u'(x"64"),u'(x"17"),u'(x"b8"),
u'(x"b8"),u'(x"10"),u'(x"b8"),u'(x"01"),u'(x"09"),u'(x"b6"),u'(x"00"),u'(x"0a"),u'(x"b8"),u'(x"09"),u'(x"b6"),u'(x"00"),u'(x"0a"),u'(x"b8"),u'(x"0a"),u'(x"0a"),
u'(x"0a"),u'(x"b8"),u'(x"8a"),u'(x"b8"),u'(x"0a"),u'(x"0a"),u'(x"15"),u'(x"b8"),u'(x"09"),u'(x"b6"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"0b"),u'(x"02"),u'(x"8a"),
u'(x"b8"),u'(x"01"),u'(x"15"),u'(x"b7"),u'(x"09"),u'(x"b0"),u'(x"86"),u'(x"0c"),u'(x"09"),u'(x"b0"),u'(x"01"),u'(x"8c"),u'(x"b8"),u'(x"86"),u'(x"0b"),u'(x"67"),
u'(x"b8"),u'(x"0c"),u'(x"00"),u'(x"47"),u'(x"0a"),u'(x"02"),u'(x"e7"),u'(x"b8"),u'(x"0c"),u'(x"1d"),u'(x"b8"),u'(x"10"),u'(x"b8"),u'(x"0a"),u'(x"03"),u'(x"01"),
u'(x"10"),u'(x"11"),u'(x"8a"),u'(x"b8"),u'(x"01"),u'(x"0b"),u'(x"03"),u'(x"11"),u'(x"b8"),u'(x"09"),u'(x"b6"),u'(x"15"),u'(x"00"),u'(x"b8"),u'(x"11"),u'(x"09"),
u'(x"b5"),u'(x"01"),u'(x"17"),u'(x"b8"),u'(x"d3"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"b8"),u'(x"01"),u'(x"0c"),u'(x"15"),u'(x"00"),u'(x"b8"),u'(x"0b"),u'(x"03"),
u'(x"11"),u'(x"b8"),u'(x"17"),u'(x"b8"),u'(x"25"),u'(x"00"),u'(x"b8"),u'(x"03"),u'(x"0c"),u'(x"87"),u'(x"1f"),u'(x"b8"),u'(x"01"),u'(x"93"),u'(x"09"),u'(x"b5"),
u'(x"01"),u'(x"09"),u'(x"b6"),u'(x"01"),u'(x"8a"),u'(x"b8"),u'(x"17"),u'(x"b8"),u'(x"03"),u'(x"09"),u'(x"b6"),u'(x"8b"),u'(x"b8"),u'(x"03"),u'(x"17"),u'(x"b8"),
u'(x"b8"),u'(x"60"),u'(x"b8"),u'(x"09"),u'(x"b6"),u'(x"17"),u'(x"b8"),u'(x"15"),u'(x"00"),u'(x"b8"),u'(x"17"),u'(x"b8"),u'(x"09"),u'(x"b5"),u'(x"13"),u'(x"b8"),
u'(x"15"),u'(x"2f"),u'(x"0a"),u'(x"03"),u'(x"00"),u'(x"09"),u'(x"b6"),u'(x"01"),u'(x"17"),u'(x"b8"),u'(x"03"),u'(x"09"),u'(x"b6"),u'(x"e0"),u'(x"b8"),u'(x"01"),
u'(x"15"),u'(x"b8"),u'(x"0c"),u'(x"0b"),u'(x"03"),u'(x"0c"),u'(x"87"),u'(x"0c"),u'(x"65"),u'(x"b8"),u'(x"0a"),u'(x"03"),u'(x"80"),u'(x"20"),u'(x"03"),u'(x"21"),
u'(x"b8"),u'(x"86"),u'(x"0b"),u'(x"01"),u'(x"11"),u'(x"01"),u'(x"0a"),u'(x"81"),u'(x"02"),u'(x"10"),u'(x"b8"),u'(x"0a"),u'(x"b8"),u'(x"01"),u'(x"0a"),u'(x"15"),
u'(x"b8"),u'(x"b8"),u'(x"15"),u'(x"b4"),u'(x"b8"),u'(x"0a"),u'(x"b8"),u'(x"0b"),u'(x"21"),u'(x"00"),u'(x"83"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"b8"),u'(x"02"),
u'(x"09"),u'(x"b6"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"e7"),u'(x"b8"),u'(x"0a"),u'(x"0a"),u'(x"11"),u'(x"09"),u'(x"b5"),u'(x"11"),u'(x"0c"),u'(x"87"),u'(x"25"),
u'(x"ff"),u'(x"06"),u'(x"25"),u'(x"00"),u'(x"05"),u'(x"0a"),u'(x"b8"),u'(x"09"),u'(x"b5"),u'(x"0a"),u'(x"b8"),u'(x"00"),u'(x"b1"),u'(x"15"),u'(x"b8"),u'(x"14"),
u'(x"14"),u'(x"12"),u'(x"20"),u'(x"82"),u'(x"00"),u'(x"0a"),u'(x"01"),u'(x"0a"),u'(x"0b"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"b8"),u'(x"17"),u'(x"b8"),u'(x"17"),
u'(x"b8"),u'(x"0a"),u'(x"20"),u'(x"b8"),u'(x"82"),u'(x"8b"),u'(x"ff"),u'(x"81"),u'(x"15"),u'(x"40"),u'(x"12"),u'(x"0b"),u'(x"02"),u'(x"41"),u'(x"41"),u'(x"20"),
u'(x"02"),u'(x"11"),u'(x"09"),u'(x"b6"),u'(x"10"),u'(x"09"),u'(x"b5"),u'(x"1d"),u'(x"00"),u'(x"09"),u'(x"b6"),u'(x"12"),u'(x"09"),u'(x"b5"),u'(x"15"),u'(x"24"),
u'(x"01"),u'(x"00"),u'(x"b1"),u'(x"09"),u'(x"b3"),u'(x"90"),u'(x"01"),u'(x"09"),u'(x"b3"),u'(x"10"),u'(x"01"),u'(x"00"),u'(x"20"),u'(x"03"),u'(x"15"),u'(x"3e"),
u'(x"10"),u'(x"0a"),u'(x"0a"),u'(x"60"),u'(x"20"),u'(x"03"),u'(x"00"),u'(x"90"),u'(x"0a"),u'(x"0c"),u'(x"60"),u'(x"20"),u'(x"01"),u'(x"0b"),u'(x"03"),u'(x"95"),
u'(x"00"),u'(x"b8"),u'(x"0c"),u'(x"87"),u'(x"0c"),u'(x"11"),u'(x"b8"),u'(x"09"),u'(x"b6"),u'(x"8a"),u'(x"b8"),u'(x"8b"),u'(x"b8"),u'(x"02"),u'(x"15"),u'(x"00"),
u'(x"1f"),u'(x"b8"),u'(x"b8"),u'(x"15"),u'(x"00"),u'(x"b8"),u'(x"0a"),u'(x"0a"),u'(x"04"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"13"),
u'(x"17"),u'(x"b8"),u'(x"45"),u'(x"00"),u'(x"93"),u'(x"ff"),u'(x"0b"),u'(x"b8"),u'(x"03"),u'(x"55"),u'(x"00"),u'(x"15"),u'(x"b4"),u'(x"00"),u'(x"15"),u'(x"00"),
u'(x"00"),u'(x"17"),u'(x"b8"),u'(x"00"),u'(x"97"),u'(x"b8"),u'(x"05"),u'(x"0b"),u'(x"02"),u'(x"0b"),u'(x"03"),u'(x"11"),u'(x"b8"),u'(x"09"),u'(x"b6"),u'(x"a7"),
u'(x"b8"),u'(x"00"),u'(x"82"),u'(x"8b"),u'(x"b8"),u'(x"02"),u'(x"8a"),u'(x"b8"),u'(x"01"),u'(x"15"),u'(x"b8"),u'(x"15"),u'(x"b8"),u'(x"95"),u'(x"00"),u'(x"b8"),
u'(x"11"),u'(x"b8"),u'(x"15"),u'(x"b8"),u'(x"11"),u'(x"11"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"97"),u'(x"b8"),u'(x"03"),u'(x"8a"),u'(x"03"),u'(x"09"),
u'(x"b6"),u'(x"00"),u'(x"8b"),u'(x"b8"),u'(x"02"),u'(x"0a"),u'(x"1d"),u'(x"b8"),u'(x"b8"),u'(x"0b"),u'(x"21"),u'(x"00"),u'(x"83"),u'(x"17"),u'(x"b8"),u'(x"8b"),
u'(x"b8"),u'(x"02"),u'(x"0b"),u'(x"11"),u'(x"b8"),u'(x"15"),u'(x"00"),u'(x"21"),u'(x"b8"),u'(x"03"),u'(x"0a"),u'(x"0a"),u'(x"04"),u'(x"09"),u'(x"b6"),u'(x"45"),
u'(x"00"),u'(x"11"),u'(x"65"),u'(x"00"),u'(x"b8"),u'(x"01"),u'(x"95"),u'(x"00"),u'(x"11"),u'(x"b8"),u'(x"91"),u'(x"b8"),u'(x"0a"),u'(x"b8"),u'(x"06"),u'(x"15"),
u'(x"00"),u'(x"b8"),u'(x"09"),u'(x"b6"),u'(x"00"),u'(x"97"),u'(x"b8"),u'(x"0c"),u'(x"65"),u'(x"3b"),u'(x"09"),u'(x"b6"),u'(x"97"),u'(x"b8"),u'(x"1d"),u'(x"b8"),
u'(x"15"),u'(x"00"),u'(x"b8"),u'(x"09"),u'(x"b5"),u'(x"00"),u'(x"b1"),u'(x"0b"),u'(x"b8"),u'(x"02"),u'(x"10"),u'(x"15"),u'(x"b8"),u'(x"15"),u'(x"b8"),u'(x"23"),
u'(x"87"),u'(x"23"),u'(x"83"),u'(x"11"),u'(x"0b"),u'(x"21"),u'(x"b8"),u'(x"87"),u'(x"e2"),u'(x"e5"),u'(x"b8"),u'(x"87"),u'(x"0c"),u'(x"65"),u'(x"2c"),u'(x"09"),
u'(x"b6"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"ff"),u'(x"25"),u'(x"00"),u'(x"b8"),u'(x"02"),u'(x"90"),u'(x"0c"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"b5"),
u'(x"09"),u'(x"b6"),u'(x"45"),u'(x"ff"),u'(x"a3"),u'(x"00"),u'(x"86"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"20"),u'(x"55"),u'(x"01"),u'(x"10"),u'(x"65"),u'(x"00"),
u'(x"0a"),u'(x"0c"),u'(x"0c"),u'(x"0a"),u'(x"02"),u'(x"65"),u'(x"20"),u'(x"09"),u'(x"b6"),u'(x"0a"),u'(x"02"),u'(x"0b"),u'(x"00"),u'(x"8b"),u'(x"ff"),u'(x"80"),
u'(x"90"),u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"0a"),u'(x"09"),u'(x"b6"),u'(x"0a"),u'(x"09"),u'(x"b6"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"01"),u'(x"8b"),u'(x"ff"),
u'(x"80"),u'(x"97"),u'(x"ff"),u'(x"00"),u'(x"09"),u'(x"b6"),u'(x"0a"),u'(x"45"),u'(x"ff"),u'(x"0a"),u'(x"03"),u'(x"a0"),u'(x"00"),u'(x"03"),u'(x"a0"),u'(x"00"),
u'(x"83"),u'(x"e5"),u'(x"00"),u'(x"09"),u'(x"b6"),u'(x"a5"),u'(x"00"),u'(x"03"),u'(x"00"),u'(x"97"),u'(x"b8"),u'(x"80"),u'(x"97"),u'(x"b8"),u'(x"01"),u'(x"8c"),
u'(x"8c"),u'(x"8c"),u'(x"8c"),u'(x"45"),u'(x"00"),u'(x"90"),u'(x"ff"),u'(x"97"),u'(x"ff"),u'(x"b8"),u'(x"97"),u'(x"ff"),u'(x"b8"),u'(x"8a"),u'(x"ff"),u'(x"8a"),
u'(x"ff"),u'(x"09"),u'(x"b6"),u'(x"95"),u'(x"03"),u'(x"09"),u'(x"b6"),u'(x"01"),u'(x"95"),u'(x"00"),u'(x"ff"),u'(x"09"),u'(x"b6"),u'(x"8b"),u'(x"ff"),u'(x"80"),
u'(x"35"),u'(x"08"),u'(x"ff"),u'(x"03"),u'(x"8b"),u'(x"ff"),u'(x"80"),u'(x"97"),u'(x"b8"),u'(x"ff"),u'(x"97"),u'(x"b8"),u'(x"ff"),u'(x"00"),u'(x"0b"),u'(x"03"),
u'(x"25"),u'(x"00"),u'(x"b8"),u'(x"03"),u'(x"82"),u'(x"11"),u'(x"b8"),u'(x"01"),u'(x"91"),u'(x"b8"),u'(x"00"),u'(x"09"),u'(x"b6"),u'(x"10"),u'(x"03"),u'(x"11"),
u'(x"02"),u'(x"17"),u'(x"b8"),u'(x"15"),u'(x"b7"),u'(x"0a"),u'(x"0a"),u'(x"09"),u'(x"0a"),u'(x"02"),u'(x"09"),u'(x"09"),u'(x"b7"),u'(x"11"),u'(x"e5"),u'(x"00"),
u'(x"09"),u'(x"b7"),u'(x"63"),u'(x"0b"),u'(x"03"),u'(x"11"),u'(x"09"),u'(x"04"),u'(x"8b"),u'(x"03"),u'(x"00"),u'(x"01"),u'(x"90"),u'(x"01"),u'(x"55"),u'(x"00"),
u'(x"ff"),u'(x"09"),u'(x"b6"),u'(x"45"),u'(x"ff"),u'(x"60"),u'(x"0a"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"09"),u'(x"00"),u'(x"50"),u'(x"00"),u'(x"0a"),u'(x"0a"),
u'(x"40"),u'(x"10"),u'(x"b8"),u'(x"09"),u'(x"8b"),u'(x"02"),u'(x"40"),u'(x"11"),u'(x"b8"),u'(x"95"),u'(x"00"),u'(x"b8"),u'(x"00"),u'(x"b1"),u'(x"09"),u'(x"b6"),
u'(x"15"),u'(x"b7"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"09"),u'(x"11"),u'(x"65"),u'(x"00"),u'(x"e1"),u'(x"09"),u'(x"11"),u'(x"09"),u'(x"21"),u'(x"86"),u'(x"95"),
u'(x"09"),u'(x"b7"),u'(x"01"),u'(x"90"),u'(x"09"),u'(x"09"),u'(x"01"),u'(x"09"),u'(x"b7"),u'(x"00"),u'(x"e0"),u'(x"00"),u'(x"b6"),u'(x"b2"),u'(x"b2"),u'(x"b0"),
u'(x"b1"),u'(x"b2"),u'(x"b2"),u'(x"b2"),u'(x"b2"),u'(x"b1"),u'(x"b1"),u'(x"b3"),u'(x"b2"),u'(x"b7"),u'(x"b3"),u'(x"b4"),u'(x"b4"),u'(x"b4"),u'(x"b6"),u'(x"b3"),
u'(x"b4"),u'(x"b0"),u'(x"b1"),u'(x"b3"),u'(x"b1"),u'(x"b2"),u'(x"b2"),u'(x"b1"),u'(x"50"),u'(x"4c"),u'(x"43"),u'(x"46"),u'(x"42"),u'(x"0a"),u'(x"21"),u'(x"2c"),
u'(x"3b"),u'(x"3e"),u'(x"42"),u'(x"44"),u'(x"46"),u'(x"49"),u'(x"4f"),u'(x"52"),u'(x"57"),u'(x"5c"),u'(x"5f"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00") 
);


begin
   base_addr_match <= '1' when base_addr(17 downto 12) = bus_addr(17 downto 12) else '0';
   bus_addr_match <= base_addr_match;

   process(clk, base_addr_match)
   begin
      if clk = '1' and clk'event then
         bus_dati(7 downto 0) <= meme(conv_integer(bus_addr(11 downto 1)));
         bus_dati(15 downto 8) <= memo(conv_integer(bus_addr(11 downto 1)));
      end if;
   end process;

   process(clk, base_addr_match)
   begin
      if clk = '1' and clk'event then
         if base_addr_match = '1' and bus_control_dato = '1' then
            if bus_control_datob = '0' or (bus_control_datob = '1' and bus_addr(0) = '0') then
               meme(conv_integer(bus_addr(11 downto 1))) <= bus_dato(7 downto 0);
            end if;
            if bus_control_datob = '0' or (bus_control_datob = '1' and bus_addr(0) = '1') then
               memo(conv_integer(bus_addr(11 downto 1))) <= bus_dato(15 downto 8);
            end if;
         end if;
      end if;
   end process;
end implementation;

