����  �  <(*!<8!2	2	> **(8!		>(*	. (8 8*. ?<-;$
*****?><(#=?+2: <;:9872	65430&2.*  228 28 2< 1> /2/o1 /  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ���@�xD��� R >r ���0��� 7� �� 7����'0�C� �0�����G��7����A� A�A��A��A� A�A��A��y� y�y���1y� y�y��y��    =  8�?�Q����$�iQ �@��!p(��q�� $^���Q�Se�R����z��F�X#$�V��R���6Ѐ5Ј���" "RP �^a�?���^����e�?$�^��?�/a?��!�?�X� ?�o���?$��凿d�Q��� ����3�<�ce�@?��@���r"  @��0��#�
 �����b��p�0���� �4 ���#�#�
0p�Tp "H�P�>@��0��� ��d�6� ? �"���w �)�l���ب/�Ѩ��9(����cށl� >��<��s!��(��d������ш�2��r��dѨ?�������2!����c����Ѥ@�@����:�8?�ѧވ����� ���&�)Ɉ  �����k �)��  0���� �� �� �� �� �� ��  ����?3 �#� �&�	&�&(?��!>�	É�Ϟ����!�		c���	�+�2 �&�J���W;����&˪'��B��s�(�����������w��'��'��'��'�����r�&|��� �� >��b� ~� ?��"�����'��KP3A�v�P3��D�T  (E� ��r��q�P�At9�GH�O8� a�                    t                      �              � p         �e	�ۀ����� �wM v�weI ��Ě�Ԡ)�Hp��窔4�x#fmU��  ���o�        �?��q����w����ty��f�� ��`�s���  ���&�'~-&'�i����/�-��<--s��� ֎ �b��x-bM�����D���C�}�*�����|��\��(��{�@����z&�������j���)`/��)Rk )���y"(��xK)L��+ 7(8�6&,�!��ԫ ��|����� ��N�|��!���/S�D�   ,P ���̀��e�-�B..g��M������ � �.�"����-�.'.�K.�"����.�-�7�/�-�~&)(/�ȯL�(��K��L~�.*f� ��,�Nz�M��!.(R�KQ�c6��x��}�������-Rk~.&-f�6�CN� ��7"���x�+�.&-fA��B��y�/-7"���B ���� .�.�.�;    � ��7Ɓ�'(/%�/���Z���#�[#��ވ�(���P5��/�5��]�����&� .&���'�hSQ�mZ�[ʖ�]��\)SO��� �� �O��� X�?'�/���Oɐ�� X'� ��Q� &��wb
vb}b�w�u9)Xv�k ��5bt�5.s�&�,r�   �޴��+ �&�,r�1  � �JKk'�/�Z����#[)#�b�&b�r�   �	]��(�� ���bb&���''b���X�?�����G@�RS�Qd�Qe�����$��'���T����R��  ��C�W��U��Qr��%��?����WϚUϚQw�u�)SO��� �%���u�)X�?'�/���{            �6�bO�k$ʦJ:k1KZ$�[$��1b�����&&�,r�   ���!�����]i��&S ����ʁ,|rq(/̛�u�+��Þك�t@��c�ك�t@J
��J.
��ӨJ���/ʎ�Ӊ��&��&��JPf���&$\)$�j   � h$�� �����O̐�(�Oϐ�� (�B�S�(Qi+ �(�/��R �,(/�!�,�k   ʼ":1�'�/�s��l�0t.����Z�%�&%�b[%�1�&2�&3�&4�&&�&����]i��&�b��b�S{%\)%Qio �       p %b����,�R�q"��϶Ը ���{�1 �
%\)%�kQ�  %�� �������K*�/�T�,�&.�&�*�S��*�/�Y��.&S*�Q��    ,�S���3��O����r��i��r��d�������t ��7�.tत7�����Z��Zu�,��{    B	�:�Y��:)�
�o�/�Ӧ���
�&v
&���l��� �`.�/��F��� /
�i��Qix �,�nNi�`/���H��	,bF,�D	�,�j�(/�������.�.,b!N� ���	Gn{B:�?T������v?S�n(/������K)�BV���"���W��U��mK)��Bw����� .�Li�J� �xK)}K)�.�,�h�&�"�?�ŉ��|W��,�Ju�,�|SP�#��.��,�0T��&�Áq�(��uC)Y(�(���Qc�UΚ E	n�/A��T�� �Nz�̨/���..&� ��k    � ��ڀ�X��,(/�,�,�/�T�BS�W��U���U��X��S� T	�R�V,�,,BȘ��,�(��,�hT.��Ni7(/�6�D��Uǒ.�j�y����R�� X	Ǻ�W���X�
"
fR �X�����ǛEǔ�E�y�/ .�+�l"���&��
�lC
t�Ϊ �	�Ƕ%!.#�/�q.�/q.ǐ/��B� ���kT� �R�� R� (��憆K߆�@����� ���EV���
l"�����F�߸�A�����R�@ ��ߨRA���R�S ��/�E�V��������R��R��S��SX����RE�k�/���,����T��RU�ה�RU�� �!.EV���K n ����� �(�n / �/�YI� �
"�l�<�Ǵ��腠���iRø�JEn������R��������!.��iRô�������R��脟E�n�/�R� ��&�&�Ni7(/��� ���t�JQ�� /�Ti� ����`/٪�
"�b�b!�(?�!��Á�����J,,B����&,�/SR� �t��N�z!��4���Qc��+�+Rk�����U  (b�'��X������a␀�
b!�@j�����(����n
&7���d��
B�z
'�
�!�PjⰀ�� ������� �
�"���F��H�� 4M�	t��&�R���b(�����ω��� �� �  H.HH��@/��iC)�J� ������r	��k   ��f���� � ���?�E�V����?�M)!����,C���M)Z�f��?��"(���@.��.�/�i�C����mC)�J�m�
��l��cV`���	fc�M�!������!.�/ڌ������k�/��w ������E�����M!��
�/���	k2���	&	7!.�/���ir� �      ^
��_� ��:��$� ����W����K ��Ͳ9��� ����W����K ���b9͒����
�o�/����hb:�����`.�/�֮&�
�l�/�� ⨩�
!.P.��/H��� ���h�/��bq�/��9͛�$�
�!�P��F�GӚ ��Á�� �
�&�
�
�l�<� �    �	 u� ���`/�������p�4t�p0�c�LtJ
��J
b|r�k�歠*�殠*      ��bH��������&���b
�
t୉,�~&�.t�'��ˁ��&���&���            ��D��D��'��'��'��'��'u�,��|����Tݟ���� �                                                                                                                                         �&~	&�Á(��|��(/��"	�z6	'	�|�<�k��'� �"#1!���� ���H/��������lp0�ctJ
���cp��<t�J
b|r�k�氤*�汤*      ��b(�����b��k���&�.tఉ,t�.

�t��|�K���&� ��
ǁ�� ��&ۉ,�|���k !��c�F(?�ࢠ���#��c��k��K �a.�/���&
	&h"�����	rh�/���I)d��&j&;�� /	�|�(�����	h"���v&	&!.
�/����<9���*P���&u9)� ��
�o�)��&g&w&!.
�/���<>i�/�w�	b!
������	�|�	�
dJ)� �q(/((/X����K� �	!.�/�
bl�/�
��hl"���I)�n&��f&j&<�(���ǁ��&�/�w�	b�j��	�|!.�/�	�
�k ��"�fbgbvb�l6�=ɠ�b���v&��!.�/���n&J)� ����|���n&� ��� ��� �   xº �v�<q�/��!!b"�h���&g&;����>�q�/�����!a.�/����/�"�!!��""BJ��P���/<u�>i� �!I)!t��j&�&�>�>"�`���""BJ��;���	�|	�"��j"���v&	&!.
�/����<9���*`.�/���nPi�Ϛ    �	��!&��"�nfbgb<i=�j�/�!�!⨵�!I)�~!!&���&b����"�""b!���"J)��f&g&��
b	bh�/���	7��� � ���4� h#��   ��� ��Xc����a.�/��a�� #��� � �����Pi R ]	�
>

�emK�emKL���KQ� 5�/&01f23f4�bdbNibM?�(��X�be��F���z1/&2�*����5�j�R� �bNizM	*�Qe� ���"�b��/4�/(?�4��Q�� �1(/�ض2�&3�&4�&��K      �,�.���(�,(/�,� ,b(S����T�@S�U�AiSU�� ��?���4�  Ɗ�{���/�&0�&�r�
     ���&�b �����&b�r�  �������+Q(� ���&��&�rB��&�(?����Q�!����&� .�������R��+ �����b�l� !�������D΁�� �   � �n��b r(/�g�gF���&��C�H?���H>(���o�߫���       | �(/��(���(/�D���&�a,���/H �C��������&��"��k��"��j ��~b�i�� ��� �d�&�c"�a,a ��J��남/�����ab�� ���,����T�c,$ւ�S �                                  @Ȁ�P���H���
�"�����&
�,�����&�l"����V9ډJ�
�!��-�/���b��x�@����!.�"(���/�ڸ�Ák�H���H/�(�+x"��������/�}��+������2�@/�!��@?����ê����֮i�*��&��� �� ���'�m�� � ,(��� ��fS��  W������D7� ̰,��E!�r��A�4��� PPfPPfPQfQQf��f��f��f��f��f��f�� ��  b�f��`�� �� �� �� �  � � #LX"2�!3�!�� �� ݛ  $(�+�.��INLEG			!�,�b,bF�,,bw��K)�JLS�                              ���/E*AU2 U][\,�/ID��USIe1K��^��N��D�� ��w�p�� �� �� �� �� �� �� �� �� �� �� �� �� �� ��  � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �  !/+�id��[�%��U�b[`���S�\E5U����"1MD �DQ4�`k3